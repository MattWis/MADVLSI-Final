magic
tech scmos
timestamp 1414783565
<< psubstratepcontact >>
rect -46 -2 -31 10
<< metal1 >>
rect -52 10 -37 47
rect -52 -1 -46 10
use Bias  Bias_0
timestamp 1414783014
transform 1 0 -262 0 1 255
box 69 -266 207 42
use FCDAmp  FCDAmp_0
timestamp 1414783254
transform 1 0 -28 0 1 92
box -27 -68 105 211
<< labels >>
rlabel metal1 -52 10 -37 47 1 Gnd
<< end >>
