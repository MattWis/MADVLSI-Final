magic
tech scmos
timestamp 1418336218
<< error_p >>
rect 182 -79 201 -22
rect 205 -79 206 -22
rect 278 -37 282 -36
rect 259 -38 261 -37
rect 267 -38 269 -37
rect 275 -38 277 -37
rect 283 -38 285 -33
rect 310 -37 314 -36
rect 291 -38 293 -37
rect 299 -38 301 -37
rect 307 -38 309 -37
rect 315 -38 317 -33
rect 323 -38 325 -37
rect 331 -38 333 -37
rect 180 -116 201 -79
rect 204 -81 206 -79
rect 180 -132 199 -116
rect 205 -126 206 -81
rect 180 -139 200 -132
rect 180 -141 205 -139
rect 180 -142 204 -141
rect 180 -151 201 -142
rect 195 -155 199 -154
rect 197 -156 199 -155
rect 197 -217 199 -216
rect 246 -217 248 -216
rect 269 -217 270 -216
rect 272 -217 273 -216
<< nwell >>
rect 189 -141 190 -79
rect 191 -116 192 -22
rect 196 -116 205 -22
rect 191 -141 205 -116
rect 189 -142 191 -141
<< polysilicon >>
rect 259 83 261 85
rect 267 83 269 85
rect 275 83 277 85
rect 283 83 285 85
rect 291 83 293 85
rect 299 83 301 85
rect 307 83 309 85
rect 315 83 317 85
rect 323 83 325 85
rect 331 83 333 85
rect 197 -21 199 -19
rect 163 -135 165 -133
rect 168 -135 170 -133
rect 178 -134 180 -132
rect 163 -149 165 -141
rect 168 -142 170 -141
rect 168 -143 174 -142
rect 168 -147 169 -143
rect 173 -147 174 -143
rect 168 -148 174 -147
rect 158 -150 165 -149
rect 158 -154 159 -150
rect 163 -154 165 -150
rect 158 -155 165 -154
rect 171 -155 174 -148
rect 178 -149 180 -146
rect 193 -147 199 -142
rect 177 -150 183 -149
rect 177 -154 178 -150
rect 182 -154 183 -150
rect 177 -155 183 -154
rect 193 -151 194 -147
rect 198 -151 199 -147
rect 193 -155 199 -151
rect 210 -143 294 -142
rect 210 -154 211 -143
rect 215 -154 294 -143
rect 210 -155 294 -154
rect 162 -156 164 -155
rect 172 -156 174 -155
rect 180 -156 182 -155
rect 214 -156 216 -155
rect 222 -156 224 -155
rect 230 -156 232 -155
rect 238 -156 240 -155
rect 246 -156 248 -155
rect 254 -156 256 -155
rect 262 -156 264 -155
rect 270 -156 272 -155
rect 278 -156 280 -155
rect 286 -156 288 -155
rect 162 -164 164 -162
rect 172 -164 174 -162
rect 180 -164 182 -162
rect 214 -218 216 -216
rect 222 -218 224 -216
rect 230 -218 232 -216
rect 238 -218 240 -216
rect 254 -218 256 -216
rect 262 -218 264 -216
rect 270 -219 272 -217
rect 278 -218 280 -216
rect 286 -218 288 -216
<< ndiffusion >>
rect 156 -157 162 -156
rect 156 -161 157 -157
rect 161 -161 162 -157
rect 156 -162 162 -161
rect 164 -157 172 -156
rect 164 -161 165 -157
rect 171 -161 172 -157
rect 164 -162 172 -161
rect 174 -157 180 -156
rect 174 -161 175 -157
rect 179 -161 180 -157
rect 174 -162 180 -161
rect 182 -157 188 -156
rect 182 -161 183 -157
rect 187 -161 188 -157
rect 182 -162 188 -161
rect 191 -157 197 -156
rect 191 -161 192 -157
rect 196 -161 197 -157
rect 165 -166 171 -162
rect 191 -165 197 -161
rect 191 -169 192 -165
rect 196 -169 197 -165
rect 191 -173 197 -169
rect 191 -177 192 -173
rect 196 -177 197 -173
rect 191 -181 197 -177
rect 191 -191 192 -181
rect 196 -191 197 -181
rect 191 -195 197 -191
rect 191 -199 192 -195
rect 196 -199 197 -195
rect 191 -203 197 -199
rect 191 -207 192 -203
rect 196 -207 197 -203
rect 191 -211 197 -207
rect 191 -215 192 -211
rect 196 -215 197 -211
rect 191 -216 197 -215
rect 199 -157 205 -156
rect 199 -215 200 -157
rect 204 -215 205 -157
rect 199 -216 205 -215
rect 208 -157 214 -156
rect 208 -161 209 -157
rect 213 -161 214 -157
rect 208 -165 214 -161
rect 208 -169 209 -165
rect 213 -169 214 -165
rect 208 -173 214 -169
rect 208 -177 209 -173
rect 213 -177 214 -173
rect 208 -181 214 -177
rect 208 -191 209 -181
rect 213 -191 214 -181
rect 208 -195 214 -191
rect 208 -199 209 -195
rect 213 -199 214 -195
rect 208 -203 214 -199
rect 208 -207 209 -203
rect 213 -207 214 -203
rect 208 -211 214 -207
rect 208 -215 209 -211
rect 213 -215 214 -211
rect 208 -216 214 -215
rect 216 -157 222 -156
rect 216 -215 217 -157
rect 221 -215 222 -157
rect 216 -216 222 -215
rect 224 -157 230 -156
rect 224 -161 225 -157
rect 229 -161 230 -157
rect 224 -165 230 -161
rect 224 -169 225 -165
rect 229 -169 230 -165
rect 224 -173 230 -169
rect 224 -177 225 -173
rect 229 -177 230 -173
rect 224 -181 230 -177
rect 224 -191 225 -181
rect 229 -191 230 -181
rect 224 -195 230 -191
rect 224 -199 225 -195
rect 229 -199 230 -195
rect 224 -203 230 -199
rect 224 -207 225 -203
rect 229 -207 230 -203
rect 224 -211 230 -207
rect 224 -215 225 -211
rect 229 -215 230 -211
rect 224 -216 230 -215
rect 232 -157 238 -156
rect 232 -215 233 -157
rect 237 -215 238 -157
rect 232 -216 238 -215
rect 240 -157 246 -156
rect 240 -161 241 -157
rect 245 -161 246 -157
rect 240 -165 246 -161
rect 240 -169 241 -165
rect 245 -169 246 -165
rect 240 -173 246 -169
rect 240 -177 241 -173
rect 245 -177 246 -173
rect 240 -181 246 -177
rect 240 -191 241 -181
rect 245 -191 246 -181
rect 240 -195 246 -191
rect 240 -199 241 -195
rect 245 -199 246 -195
rect 240 -203 246 -199
rect 240 -207 241 -203
rect 245 -207 246 -203
rect 240 -211 246 -207
rect 240 -215 241 -211
rect 245 -215 246 -211
rect 240 -216 246 -215
rect 248 -157 254 -156
rect 248 -215 249 -157
rect 253 -215 254 -157
rect 248 -216 254 -215
rect 256 -157 262 -156
rect 256 -161 257 -157
rect 261 -161 262 -157
rect 256 -165 262 -161
rect 256 -169 257 -165
rect 261 -169 262 -165
rect 256 -173 262 -169
rect 256 -177 257 -173
rect 261 -177 262 -173
rect 256 -181 262 -177
rect 256 -191 257 -181
rect 261 -191 262 -181
rect 256 -195 262 -191
rect 256 -199 257 -195
rect 261 -199 262 -195
rect 256 -203 262 -199
rect 256 -207 257 -203
rect 261 -207 262 -203
rect 256 -211 262 -207
rect 256 -215 257 -211
rect 261 -215 262 -211
rect 256 -216 262 -215
rect 264 -157 270 -156
rect 264 -215 265 -157
rect 269 -215 270 -157
rect 264 -216 270 -215
rect 272 -157 278 -156
rect 272 -161 273 -157
rect 277 -161 278 -157
rect 272 -165 278 -161
rect 272 -169 273 -165
rect 277 -169 278 -165
rect 272 -173 278 -169
rect 272 -177 273 -173
rect 277 -177 278 -173
rect 272 -181 278 -177
rect 272 -191 273 -181
rect 277 -191 278 -181
rect 272 -195 278 -191
rect 272 -199 273 -195
rect 277 -199 278 -195
rect 272 -203 278 -199
rect 272 -207 273 -203
rect 277 -207 278 -203
rect 272 -211 278 -207
rect 272 -215 273 -211
rect 277 -215 278 -211
rect 272 -216 278 -215
rect 280 -157 286 -156
rect 280 -215 281 -157
rect 285 -215 286 -157
rect 280 -216 286 -215
rect 288 -157 294 -156
rect 288 -161 289 -157
rect 293 -161 294 -157
rect 288 -165 294 -161
rect 288 -169 289 -165
rect 293 -169 294 -165
rect 288 -173 294 -169
rect 288 -177 289 -173
rect 293 -177 294 -173
rect 288 -181 294 -177
rect 288 -191 289 -181
rect 293 -191 294 -181
rect 288 -195 294 -191
rect 288 -199 289 -195
rect 293 -199 294 -195
rect 288 -203 294 -199
rect 288 -207 289 -203
rect 293 -207 294 -203
rect 288 -211 294 -207
rect 288 -215 289 -211
rect 293 -215 294 -211
rect 288 -216 294 -215
<< pdiffusion >>
rect 253 82 259 83
rect 253 76 254 82
rect 258 76 259 82
rect 253 72 259 76
rect 253 68 254 72
rect 258 68 259 72
rect 253 64 259 68
rect 253 60 254 64
rect 258 60 259 64
rect 253 56 259 60
rect 253 52 254 56
rect 258 52 259 56
rect 253 48 259 52
rect 253 44 254 48
rect 258 44 259 48
rect 253 40 259 44
rect 253 36 254 40
rect 258 36 259 40
rect 253 32 259 36
rect 253 28 254 32
rect 258 28 259 32
rect 253 24 259 28
rect 253 20 254 24
rect 258 20 259 24
rect 253 16 259 20
rect 253 12 254 16
rect 258 12 259 16
rect 253 8 259 12
rect 253 4 254 8
rect 258 4 259 8
rect 253 0 259 4
rect 253 -4 254 0
rect 258 -4 259 0
rect 253 -8 259 -4
rect 253 -12 254 -8
rect 258 -12 259 -8
rect 253 -16 259 -12
rect 253 -20 254 -16
rect 258 -20 259 -16
rect 191 -24 197 -21
rect 191 -28 192 -24
rect 196 -28 197 -24
rect 191 -32 197 -28
rect 191 -36 192 -32
rect 196 -36 197 -32
rect 191 -40 197 -36
rect 191 -44 192 -40
rect 196 -44 197 -40
rect 191 -48 197 -44
rect 191 -52 192 -48
rect 196 -52 197 -48
rect 191 -56 197 -52
rect 191 -60 192 -56
rect 196 -60 197 -56
rect 191 -64 197 -60
rect 191 -68 192 -64
rect 196 -68 197 -64
rect 191 -72 197 -68
rect 191 -76 192 -72
rect 196 -76 197 -72
rect 191 -80 197 -76
rect 191 -84 192 -80
rect 196 -84 197 -80
rect 191 -88 197 -84
rect 191 -92 192 -88
rect 196 -92 197 -88
rect 191 -96 197 -92
rect 191 -100 192 -96
rect 196 -100 197 -96
rect 191 -104 197 -100
rect 191 -108 192 -104
rect 196 -108 197 -104
rect 191 -112 197 -108
rect 191 -116 192 -112
rect 196 -116 197 -112
rect 191 -120 197 -116
rect 191 -124 192 -120
rect 196 -124 197 -120
rect 191 -128 197 -124
rect 191 -132 192 -128
rect 196 -132 197 -128
rect 175 -135 178 -134
rect 153 -136 163 -135
rect 153 -140 158 -136
rect 162 -140 163 -136
rect 153 -141 163 -140
rect 165 -141 168 -135
rect 170 -136 178 -135
rect 170 -140 172 -136
rect 176 -140 178 -136
rect 170 -141 178 -140
rect 175 -146 178 -141
rect 180 -136 186 -134
rect 180 -140 181 -136
rect 185 -140 186 -136
rect 180 -146 186 -140
rect 191 -136 197 -132
rect 191 -140 192 -136
rect 196 -140 197 -136
rect 191 -141 197 -140
rect 199 -22 205 -21
rect 199 -140 200 -22
rect 204 -140 205 -22
rect 253 -24 259 -20
rect 253 -28 254 -24
rect 258 -28 259 -24
rect 253 -32 259 -28
rect 253 -36 254 -32
rect 258 -36 259 -32
rect 253 -37 259 -36
rect 261 82 267 83
rect 261 -36 262 82
rect 266 -36 267 82
rect 261 -37 267 -36
rect 269 82 275 83
rect 269 76 270 82
rect 274 76 275 82
rect 269 72 275 76
rect 269 68 270 72
rect 274 68 275 72
rect 269 64 275 68
rect 269 60 270 64
rect 274 60 275 64
rect 269 56 275 60
rect 269 52 270 56
rect 274 52 275 56
rect 269 48 275 52
rect 269 44 270 48
rect 274 44 275 48
rect 269 40 275 44
rect 269 36 270 40
rect 274 36 275 40
rect 269 32 275 36
rect 269 28 270 32
rect 274 28 275 32
rect 269 24 275 28
rect 269 20 270 24
rect 274 20 275 24
rect 269 16 275 20
rect 269 12 270 16
rect 274 12 275 16
rect 269 8 275 12
rect 269 4 270 8
rect 274 4 275 8
rect 269 0 275 4
rect 269 -4 270 0
rect 274 -4 275 0
rect 269 -8 275 -4
rect 269 -12 270 -8
rect 274 -12 275 -8
rect 269 -16 275 -12
rect 269 -20 270 -16
rect 274 -20 275 -16
rect 269 -24 275 -20
rect 269 -28 270 -24
rect 274 -28 275 -24
rect 269 -32 275 -28
rect 269 -36 270 -32
rect 274 -36 275 -32
rect 269 -37 275 -36
rect 277 82 283 83
rect 277 -37 278 82
rect 282 -37 283 82
rect 285 82 291 83
rect 285 76 286 82
rect 290 76 291 82
rect 285 72 291 76
rect 285 68 286 72
rect 290 68 291 72
rect 285 64 291 68
rect 285 60 286 64
rect 290 60 291 64
rect 285 56 291 60
rect 285 52 286 56
rect 290 52 291 56
rect 285 48 291 52
rect 285 44 286 48
rect 290 44 291 48
rect 285 40 291 44
rect 285 36 286 40
rect 290 36 291 40
rect 285 32 291 36
rect 285 28 286 32
rect 290 28 291 32
rect 285 24 291 28
rect 285 20 286 24
rect 290 20 291 24
rect 285 16 291 20
rect 285 12 286 16
rect 290 12 291 16
rect 285 8 291 12
rect 285 4 286 8
rect 290 4 291 8
rect 285 0 291 4
rect 285 -4 286 0
rect 290 -4 291 0
rect 285 -8 291 -4
rect 285 -12 286 -8
rect 290 -12 291 -8
rect 285 -16 291 -12
rect 285 -20 286 -16
rect 290 -20 291 -16
rect 285 -24 291 -20
rect 285 -28 286 -24
rect 290 -28 291 -24
rect 285 -32 291 -28
rect 285 -36 286 -32
rect 290 -36 291 -32
rect 285 -37 291 -36
rect 293 82 299 83
rect 293 -36 294 82
rect 298 -36 299 82
rect 293 -37 299 -36
rect 301 82 307 83
rect 301 76 302 82
rect 306 76 307 82
rect 301 72 307 76
rect 301 68 302 72
rect 306 68 307 72
rect 301 64 307 68
rect 301 60 302 64
rect 306 60 307 64
rect 301 56 307 60
rect 301 52 302 56
rect 306 52 307 56
rect 301 48 307 52
rect 301 44 302 48
rect 306 44 307 48
rect 301 40 307 44
rect 301 36 302 40
rect 306 36 307 40
rect 301 32 307 36
rect 301 28 302 32
rect 306 28 307 32
rect 301 24 307 28
rect 301 20 302 24
rect 306 20 307 24
rect 301 16 307 20
rect 301 12 302 16
rect 306 12 307 16
rect 301 8 307 12
rect 301 4 302 8
rect 306 4 307 8
rect 301 0 307 4
rect 301 -4 302 0
rect 306 -4 307 0
rect 301 -8 307 -4
rect 301 -12 302 -8
rect 306 -12 307 -8
rect 301 -16 307 -12
rect 301 -20 302 -16
rect 306 -20 307 -16
rect 301 -24 307 -20
rect 301 -28 302 -24
rect 306 -28 307 -24
rect 301 -32 307 -28
rect 301 -36 302 -32
rect 306 -36 307 -32
rect 301 -37 307 -36
rect 309 82 315 83
rect 309 -37 310 82
rect 314 -37 315 82
rect 317 82 323 83
rect 317 76 318 82
rect 322 76 323 82
rect 317 72 323 76
rect 317 68 318 72
rect 322 68 323 72
rect 317 64 323 68
rect 317 60 318 64
rect 322 60 323 64
rect 317 56 323 60
rect 317 52 318 56
rect 322 52 323 56
rect 317 48 323 52
rect 317 44 318 48
rect 322 44 323 48
rect 317 40 323 44
rect 317 36 318 40
rect 322 36 323 40
rect 317 32 323 36
rect 317 28 318 32
rect 322 28 323 32
rect 317 24 323 28
rect 317 20 318 24
rect 322 20 323 24
rect 317 16 323 20
rect 317 12 318 16
rect 322 12 323 16
rect 317 8 323 12
rect 317 4 318 8
rect 322 4 323 8
rect 317 0 323 4
rect 317 -4 318 0
rect 322 -4 323 0
rect 317 -8 323 -4
rect 317 -12 318 -8
rect 322 -12 323 -8
rect 317 -16 323 -12
rect 317 -20 318 -16
rect 322 -20 323 -16
rect 317 -24 323 -20
rect 317 -28 318 -24
rect 322 -28 323 -24
rect 317 -32 323 -28
rect 317 -36 318 -32
rect 322 -36 323 -32
rect 317 -37 323 -36
rect 325 82 331 83
rect 325 -36 326 82
rect 330 -36 331 82
rect 325 -37 331 -36
rect 333 82 339 83
rect 333 76 334 82
rect 338 76 339 82
rect 333 72 339 76
rect 333 68 334 72
rect 338 68 339 72
rect 333 64 339 68
rect 333 60 334 64
rect 338 60 339 64
rect 333 56 339 60
rect 333 52 334 56
rect 338 52 339 56
rect 333 48 339 52
rect 333 44 334 48
rect 338 44 339 48
rect 333 40 339 44
rect 333 36 334 40
rect 338 36 339 40
rect 333 32 339 36
rect 333 28 334 32
rect 338 28 339 32
rect 333 24 339 28
rect 333 20 334 24
rect 338 20 339 24
rect 333 16 339 20
rect 333 12 334 16
rect 338 12 339 16
rect 333 8 339 12
rect 333 4 334 8
rect 338 4 339 8
rect 333 0 339 4
rect 333 -4 334 0
rect 338 -4 339 0
rect 333 -8 339 -4
rect 333 -12 334 -8
rect 338 -12 339 -8
rect 333 -16 339 -12
rect 333 -20 334 -16
rect 338 -20 339 -16
rect 333 -24 339 -20
rect 333 -28 334 -24
rect 338 -28 339 -24
rect 333 -32 339 -28
rect 333 -36 334 -32
rect 338 -36 339 -32
rect 333 -37 339 -36
rect 199 -141 205 -140
<< metal1 >>
rect 191 -73 192 -22
rect 150 -83 190 -82
rect 150 -130 162 -83
rect 150 -133 190 -130
rect 191 -133 192 -82
rect 170 -136 178 -133
rect 170 -140 172 -136
rect 176 -140 178 -136
rect 150 -147 169 -143
rect 185 -147 189 -136
rect 204 -81 205 -22
rect 253 -36 254 82
rect 266 -36 267 82
rect 262 -37 267 -36
rect 282 -37 283 82
rect 298 -36 299 82
rect 294 -37 299 -36
rect 314 -37 315 82
rect 330 -36 331 82
rect 326 -37 331 -36
rect 204 -140 205 -82
rect 200 -141 205 -140
rect 200 -143 205 -142
rect 218 -143 222 -142
rect 234 -143 238 -142
rect 250 -143 254 -142
rect 266 -143 270 -142
rect 282 -143 286 -142
rect 200 -144 211 -143
rect 150 -154 159 -150
rect 166 -154 178 -150
rect 185 -151 194 -147
rect 166 -157 170 -154
rect 185 -157 189 -151
rect 201 -154 211 -144
rect 218 -154 300 -143
rect 200 -157 205 -154
rect 218 -157 222 -154
rect 234 -157 238 -154
rect 250 -157 254 -154
rect 266 -157 270 -154
rect 282 -157 286 -154
rect 150 -161 157 -157
rect 187 -161 189 -157
rect 150 -169 161 -161
rect 175 -169 179 -161
rect 150 -170 192 -169
rect 150 -216 151 -170
rect 191 -215 192 -170
rect 204 -215 205 -157
rect 221 -215 222 -157
rect 237 -215 238 -157
rect 253 -215 254 -157
rect 269 -215 270 -157
rect 285 -215 286 -157
rect 191 -216 196 -215
rect 150 -217 196 -216
<< metal2 >>
rect 253 76 345 82
rect 253 72 254 76
rect 258 72 270 76
rect 274 72 286 76
rect 290 72 302 76
rect 306 72 318 76
rect 322 72 334 76
rect 338 72 345 76
rect 253 68 345 72
rect 253 64 254 68
rect 258 64 270 68
rect 274 64 286 68
rect 290 64 302 68
rect 306 64 318 68
rect 322 64 334 68
rect 338 64 345 68
rect 253 60 345 64
rect 253 56 254 60
rect 258 56 270 60
rect 274 56 286 60
rect 290 56 302 60
rect 306 56 318 60
rect 322 56 334 60
rect 338 56 345 60
rect 253 52 345 56
rect 253 48 254 52
rect 258 48 270 52
rect 274 48 286 52
rect 290 48 302 52
rect 306 48 318 52
rect 322 48 334 52
rect 338 48 345 52
rect 253 44 345 48
rect 253 40 254 44
rect 258 40 270 44
rect 274 40 286 44
rect 290 40 302 44
rect 306 40 318 44
rect 322 40 334 44
rect 338 40 345 44
rect 253 36 345 40
rect 253 32 254 36
rect 258 32 270 36
rect 274 32 286 36
rect 290 32 302 36
rect 306 32 318 36
rect 322 32 334 36
rect 338 32 345 36
rect 253 28 345 32
rect 253 24 254 28
rect 258 24 270 28
rect 274 24 286 28
rect 290 24 302 28
rect 306 24 318 28
rect 322 24 334 28
rect 338 24 345 28
rect 253 20 345 24
rect 253 16 254 20
rect 258 16 270 20
rect 274 16 286 20
rect 290 16 302 20
rect 306 16 318 20
rect 322 16 334 20
rect 338 16 345 20
rect 253 12 345 16
rect 253 8 254 12
rect 258 8 270 12
rect 274 8 286 12
rect 290 8 302 12
rect 306 8 318 12
rect 322 8 334 12
rect 338 8 345 12
rect 253 4 345 8
rect 253 0 254 4
rect 258 0 270 4
rect 274 0 286 4
rect 290 0 302 4
rect 306 0 318 4
rect 322 0 334 4
rect 338 0 345 4
rect 253 -4 345 0
rect 253 -8 254 -4
rect 258 -8 270 -4
rect 274 -8 286 -4
rect 290 -8 302 -4
rect 306 -8 318 -4
rect 322 -8 334 -4
rect 338 -8 345 -4
rect 253 -12 345 -8
rect 253 -16 254 -12
rect 258 -16 270 -12
rect 274 -16 286 -12
rect 290 -16 302 -12
rect 306 -16 318 -12
rect 322 -16 334 -12
rect 338 -16 345 -12
rect 253 -20 345 -16
rect 192 -28 205 -22
rect 196 -32 205 -28
rect 192 -36 205 -32
rect 253 -24 254 -20
rect 258 -24 270 -20
rect 274 -24 286 -20
rect 290 -24 302 -20
rect 306 -24 318 -20
rect 322 -24 334 -20
rect 338 -24 345 -20
rect 253 -28 345 -24
rect 253 -32 254 -28
rect 258 -32 270 -28
rect 274 -32 286 -28
rect 290 -32 302 -28
rect 306 -32 318 -28
rect 322 -32 334 -28
rect 338 -32 345 -28
rect 253 -36 345 -32
rect 196 -40 205 -36
rect 192 -44 205 -40
rect 196 -48 205 -44
rect 192 -52 205 -48
rect 196 -56 205 -52
rect 192 -60 205 -56
rect 196 -64 205 -60
rect 192 -68 205 -64
rect 196 -72 205 -68
rect 192 -76 205 -72
rect 196 -80 205 -76
rect 192 -84 205 -80
rect 196 -88 205 -84
rect 192 -92 205 -88
rect 196 -96 205 -92
rect 192 -100 205 -96
rect 196 -104 205 -100
rect 192 -108 205 -104
rect 196 -112 205 -108
rect 192 -116 205 -112
rect 196 -120 205 -116
rect 192 -124 205 -120
rect 196 -128 205 -124
rect 192 -132 205 -128
rect 196 -136 205 -132
rect 158 -147 162 -136
rect 192 -140 205 -136
rect 158 -151 170 -147
rect 166 -157 170 -151
rect 165 -161 170 -157
rect 192 -161 293 -157
rect 196 -165 209 -161
rect 213 -165 225 -161
rect 229 -165 241 -161
rect 245 -165 257 -161
rect 261 -165 273 -161
rect 277 -165 289 -161
rect 192 -169 293 -165
rect 196 -173 209 -169
rect 213 -173 225 -169
rect 229 -173 241 -169
rect 245 -173 257 -169
rect 261 -173 273 -169
rect 277 -173 289 -169
rect 192 -177 293 -173
rect 196 -181 209 -177
rect 213 -181 225 -177
rect 229 -181 241 -177
rect 245 -181 257 -177
rect 261 -181 273 -177
rect 277 -181 289 -177
rect 192 -191 293 -181
rect 196 -195 209 -191
rect 213 -195 225 -191
rect 229 -195 241 -191
rect 245 -195 257 -191
rect 261 -195 273 -191
rect 277 -195 289 -191
rect 192 -199 293 -195
rect 196 -203 209 -199
rect 213 -203 225 -199
rect 229 -203 241 -199
rect 245 -203 257 -199
rect 261 -203 273 -199
rect 277 -203 289 -199
rect 192 -207 293 -203
rect 196 -211 209 -207
rect 213 -211 225 -207
rect 229 -211 241 -207
rect 245 -211 257 -207
rect 261 -211 273 -207
rect 277 -211 289 -207
rect 192 -215 293 -211
<< ntransistor >>
rect 162 -162 164 -156
rect 172 -162 174 -156
rect 180 -162 182 -156
rect 197 -216 199 -156
rect 214 -216 216 -156
rect 222 -216 224 -156
rect 230 -216 232 -156
rect 238 -216 240 -156
rect 246 -216 248 -156
rect 254 -216 256 -156
rect 262 -216 264 -156
rect 270 -217 272 -156
rect 278 -216 280 -156
rect 286 -216 288 -156
<< ptransistor >>
rect 163 -141 165 -135
rect 168 -141 170 -135
rect 178 -146 180 -134
rect 197 -141 199 -21
rect 259 -37 261 83
rect 267 -37 269 83
rect 275 -37 277 83
rect 283 -37 285 83
rect 291 -37 293 83
rect 299 -37 301 83
rect 307 -37 309 83
rect 315 -37 317 83
rect 323 -37 325 83
rect 331 -37 333 83
<< polycontact >>
rect 169 -147 173 -143
rect 159 -154 163 -150
rect 178 -154 182 -150
rect 194 -151 198 -147
rect 211 -154 215 -143
<< ndcontact >>
rect 157 -161 161 -157
rect 165 -161 171 -157
rect 175 -161 179 -157
rect 183 -161 187 -157
rect 192 -161 196 -157
rect 192 -169 196 -165
rect 192 -177 196 -173
rect 192 -191 196 -181
rect 192 -199 196 -195
rect 192 -207 196 -203
rect 192 -215 196 -211
rect 200 -215 204 -157
rect 209 -161 213 -157
rect 209 -169 213 -165
rect 209 -177 213 -173
rect 209 -191 213 -181
rect 209 -199 213 -195
rect 209 -207 213 -203
rect 209 -215 213 -211
rect 217 -215 221 -157
rect 225 -161 229 -157
rect 225 -169 229 -165
rect 225 -177 229 -173
rect 225 -191 229 -181
rect 225 -199 229 -195
rect 225 -207 229 -203
rect 225 -215 229 -211
rect 233 -215 237 -157
rect 241 -161 245 -157
rect 241 -169 245 -165
rect 241 -177 245 -173
rect 241 -191 245 -181
rect 241 -199 245 -195
rect 241 -207 245 -203
rect 241 -215 245 -211
rect 249 -215 253 -157
rect 257 -161 261 -157
rect 257 -169 261 -165
rect 257 -177 261 -173
rect 257 -191 261 -181
rect 257 -199 261 -195
rect 257 -207 261 -203
rect 257 -215 261 -211
rect 265 -215 269 -157
rect 273 -161 277 -157
rect 273 -169 277 -165
rect 273 -177 277 -173
rect 273 -191 277 -181
rect 273 -199 277 -195
rect 273 -207 277 -203
rect 273 -215 277 -211
rect 281 -215 285 -157
rect 289 -161 293 -157
rect 289 -169 293 -165
rect 289 -177 293 -173
rect 289 -191 293 -181
rect 289 -199 293 -195
rect 289 -207 293 -203
rect 289 -215 293 -211
<< pdcontact >>
rect 254 76 258 82
rect 254 68 258 72
rect 254 60 258 64
rect 254 52 258 56
rect 254 44 258 48
rect 254 36 258 40
rect 254 28 258 32
rect 254 20 258 24
rect 254 12 258 16
rect 254 4 258 8
rect 254 -4 258 0
rect 254 -12 258 -8
rect 254 -20 258 -16
rect 192 -28 196 -24
rect 192 -36 196 -32
rect 192 -44 196 -40
rect 192 -52 196 -48
rect 192 -60 196 -56
rect 192 -68 196 -64
rect 192 -76 196 -72
rect 192 -84 196 -80
rect 192 -92 196 -88
rect 192 -100 196 -96
rect 192 -108 196 -104
rect 192 -116 196 -112
rect 192 -124 196 -120
rect 192 -132 196 -128
rect 158 -140 162 -136
rect 172 -140 176 -136
rect 181 -140 185 -136
rect 192 -140 196 -136
rect 200 -140 204 -22
rect 254 -28 258 -24
rect 254 -36 258 -32
rect 262 -36 266 82
rect 270 76 274 82
rect 270 68 274 72
rect 270 60 274 64
rect 270 52 274 56
rect 270 44 274 48
rect 270 36 274 40
rect 270 28 274 32
rect 270 20 274 24
rect 270 12 274 16
rect 270 4 274 8
rect 270 -4 274 0
rect 270 -12 274 -8
rect 270 -20 274 -16
rect 270 -28 274 -24
rect 270 -36 274 -32
rect 278 -36 282 82
rect 286 76 290 82
rect 286 68 290 72
rect 286 60 290 64
rect 286 52 290 56
rect 286 44 290 48
rect 286 36 290 40
rect 286 28 290 32
rect 286 20 290 24
rect 286 12 290 16
rect 286 4 290 8
rect 286 -4 290 0
rect 286 -12 290 -8
rect 286 -20 290 -16
rect 286 -28 290 -24
rect 286 -36 290 -32
rect 294 -36 298 82
rect 302 76 306 82
rect 302 68 306 72
rect 302 60 306 64
rect 302 52 306 56
rect 302 44 306 48
rect 302 36 306 40
rect 302 28 306 32
rect 302 20 306 24
rect 302 12 306 16
rect 302 4 306 8
rect 302 -4 306 0
rect 302 -12 306 -8
rect 302 -20 306 -16
rect 302 -28 306 -24
rect 302 -36 306 -32
rect 310 -36 314 82
rect 318 76 322 82
rect 318 68 322 72
rect 318 60 322 64
rect 318 52 322 56
rect 318 44 322 48
rect 318 36 322 40
rect 318 28 322 32
rect 318 20 322 24
rect 318 12 322 16
rect 318 4 322 8
rect 318 -4 322 0
rect 318 -12 322 -8
rect 318 -20 322 -16
rect 318 -28 322 -24
rect 318 -36 322 -32
rect 326 -36 330 82
rect 334 76 338 82
rect 334 68 338 72
rect 334 60 338 64
rect 334 52 338 56
rect 334 44 338 48
rect 334 36 338 40
rect 334 28 338 32
rect 334 20 338 24
rect 334 12 338 16
rect 334 4 338 8
rect 334 -4 338 0
rect 334 -12 338 -8
rect 334 -20 338 -16
rect 334 -28 338 -24
rect 334 -36 338 -32
<< m2contact >>
rect 192 -32 196 -28
rect 192 -40 196 -36
rect 192 -48 196 -44
rect 192 -56 196 -52
rect 192 -64 196 -60
rect 192 -72 196 -68
rect 192 -80 196 -76
rect 192 -88 196 -84
rect 192 -96 196 -92
rect 192 -104 196 -100
rect 192 -112 196 -108
rect 192 -120 196 -116
rect 192 -128 196 -124
rect 192 -136 196 -132
rect 154 -140 158 -136
rect 254 72 258 76
rect 254 64 258 68
rect 254 56 258 60
rect 254 48 258 52
rect 254 40 258 44
rect 254 32 258 36
rect 254 24 258 28
rect 254 16 258 20
rect 254 8 258 12
rect 254 0 258 4
rect 254 -8 258 -4
rect 254 -16 258 -12
rect 254 -24 258 -20
rect 254 -32 258 -28
rect 270 72 274 76
rect 270 64 274 68
rect 270 56 274 60
rect 270 48 274 52
rect 270 40 274 44
rect 270 32 274 36
rect 270 24 274 28
rect 270 16 274 20
rect 270 8 274 12
rect 270 0 274 4
rect 270 -8 274 -4
rect 270 -16 274 -12
rect 270 -24 274 -20
rect 270 -32 274 -28
rect 286 72 290 76
rect 286 64 290 68
rect 286 56 290 60
rect 286 48 290 52
rect 286 40 290 44
rect 286 32 290 36
rect 286 24 290 28
rect 286 16 290 20
rect 286 8 290 12
rect 286 0 290 4
rect 286 -8 290 -4
rect 286 -16 290 -12
rect 286 -24 290 -20
rect 286 -32 290 -28
rect 302 72 306 76
rect 302 64 306 68
rect 302 56 306 60
rect 302 48 306 52
rect 302 40 306 44
rect 302 32 306 36
rect 302 24 306 28
rect 302 16 306 20
rect 302 8 306 12
rect 302 0 306 4
rect 302 -8 306 -4
rect 302 -16 306 -12
rect 302 -24 306 -20
rect 302 -32 306 -28
rect 318 72 322 76
rect 318 64 322 68
rect 318 56 322 60
rect 318 48 322 52
rect 318 40 322 44
rect 318 32 322 36
rect 318 24 322 28
rect 318 16 322 20
rect 318 8 322 12
rect 318 0 322 4
rect 318 -8 322 -4
rect 318 -16 322 -12
rect 318 -24 322 -20
rect 318 -32 322 -28
rect 334 72 338 76
rect 334 64 338 68
rect 334 56 338 60
rect 334 48 338 52
rect 334 40 338 44
rect 334 32 338 36
rect 334 24 338 28
rect 334 16 338 20
rect 334 8 338 12
rect 334 0 338 4
rect 334 -8 338 -4
rect 334 -16 338 -12
rect 334 -24 338 -20
rect 334 -32 338 -28
rect 166 -165 170 -161
rect 192 -165 196 -161
rect 192 -173 196 -169
rect 192 -181 196 -177
rect 192 -195 196 -191
rect 192 -203 196 -199
rect 192 -211 196 -207
rect 209 -165 213 -161
rect 209 -173 213 -169
rect 209 -181 213 -177
rect 209 -195 213 -191
rect 209 -203 213 -199
rect 209 -211 213 -207
rect 225 -165 229 -161
rect 225 -173 229 -169
rect 225 -181 229 -177
rect 225 -195 229 -191
rect 225 -203 229 -199
rect 225 -211 229 -207
rect 241 -165 245 -161
rect 241 -173 245 -169
rect 241 -181 245 -177
rect 241 -195 245 -191
rect 241 -203 245 -199
rect 241 -211 245 -207
rect 257 -165 261 -161
rect 257 -173 261 -169
rect 257 -181 261 -177
rect 257 -195 261 -191
rect 257 -203 261 -199
rect 257 -211 261 -207
rect 273 -165 277 -161
rect 273 -173 277 -169
rect 273 -181 277 -177
rect 273 -195 277 -191
rect 273 -203 277 -199
rect 273 -211 277 -207
rect 289 -165 293 -161
rect 289 -173 293 -169
rect 289 -181 293 -177
rect 289 -195 293 -191
rect 289 -203 293 -199
rect 289 -211 293 -207
<< psubstratepcontact >>
rect 151 -216 191 -170
<< nsubstratencontact >>
rect 162 -130 190 -83
<< labels >>
rlabel metal1 155 -154 159 -150 1 B
rlabel metal1 155 -147 169 -143 1 A
rlabel metal1 218 -154 300 -143 1 Z
rlabel metal1 154 -161 157 -157 1 Gnd
<< end >>
