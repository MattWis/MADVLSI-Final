magic
tech scmos
timestamp 1418826157
<< nwell >>
rect 3370 4228 3515 4378
<< ptransistor >>
rect 3398 4245 3404 4365
rect 3419 4245 3425 4365
rect 3440 4245 3446 4365
<< pdiffusion >>
rect 3392 4364 3398 4365
rect 3392 4290 3393 4364
rect 3397 4290 3398 4364
rect 3392 4268 3398 4290
rect 3392 4246 3393 4268
rect 3397 4246 3398 4268
rect 3392 4245 3398 4246
rect 3404 4364 3410 4365
rect 3404 4358 3405 4364
rect 3409 4358 3410 4364
rect 3404 4354 3410 4358
rect 3404 4350 3405 4354
rect 3409 4350 3410 4354
rect 3404 4346 3410 4350
rect 3404 4342 3405 4346
rect 3409 4342 3410 4346
rect 3404 4338 3410 4342
rect 3404 4334 3405 4338
rect 3409 4334 3410 4338
rect 3404 4330 3410 4334
rect 3404 4326 3405 4330
rect 3409 4326 3410 4330
rect 3404 4322 3410 4326
rect 3404 4318 3405 4322
rect 3409 4318 3410 4322
rect 3404 4314 3410 4318
rect 3404 4310 3405 4314
rect 3409 4310 3410 4314
rect 3404 4306 3410 4310
rect 3404 4302 3405 4306
rect 3409 4302 3410 4306
rect 3404 4298 3410 4302
rect 3404 4294 3405 4298
rect 3409 4294 3410 4298
rect 3404 4290 3410 4294
rect 3404 4286 3405 4290
rect 3409 4286 3410 4290
rect 3404 4282 3410 4286
rect 3404 4278 3405 4282
rect 3409 4278 3410 4282
rect 3404 4274 3410 4278
rect 3404 4270 3405 4274
rect 3409 4270 3410 4274
rect 3404 4266 3410 4270
rect 3404 4262 3405 4266
rect 3409 4262 3410 4266
rect 3404 4258 3410 4262
rect 3404 4254 3405 4258
rect 3409 4254 3410 4258
rect 3404 4250 3410 4254
rect 3404 4246 3405 4250
rect 3409 4246 3410 4250
rect 3404 4245 3410 4246
rect 3413 4364 3419 4365
rect 3413 4246 3414 4364
rect 3418 4246 3419 4364
rect 3413 4245 3419 4246
rect 3425 4364 3431 4365
rect 3425 4358 3426 4364
rect 3430 4358 3431 4364
rect 3425 4354 3431 4358
rect 3425 4350 3426 4354
rect 3430 4350 3431 4354
rect 3425 4346 3431 4350
rect 3425 4342 3426 4346
rect 3430 4342 3431 4346
rect 3425 4338 3431 4342
rect 3425 4334 3426 4338
rect 3430 4334 3431 4338
rect 3425 4330 3431 4334
rect 3425 4326 3426 4330
rect 3430 4326 3431 4330
rect 3425 4322 3431 4326
rect 3425 4318 3426 4322
rect 3430 4318 3431 4322
rect 3425 4314 3431 4318
rect 3425 4310 3426 4314
rect 3430 4310 3431 4314
rect 3425 4306 3431 4310
rect 3425 4302 3426 4306
rect 3430 4302 3431 4306
rect 3425 4298 3431 4302
rect 3425 4294 3426 4298
rect 3430 4294 3431 4298
rect 3425 4290 3431 4294
rect 3425 4286 3426 4290
rect 3430 4286 3431 4290
rect 3425 4282 3431 4286
rect 3425 4278 3426 4282
rect 3430 4278 3431 4282
rect 3425 4274 3431 4278
rect 3425 4270 3426 4274
rect 3430 4270 3431 4274
rect 3425 4266 3431 4270
rect 3425 4262 3426 4266
rect 3430 4262 3431 4266
rect 3425 4258 3431 4262
rect 3425 4254 3426 4258
rect 3430 4254 3431 4258
rect 3425 4250 3431 4254
rect 3425 4246 3426 4250
rect 3430 4246 3431 4250
rect 3425 4245 3431 4246
rect 3434 4364 3440 4365
rect 3434 4246 3435 4364
rect 3439 4246 3440 4364
rect 3434 4245 3440 4246
rect 3446 4364 3452 4365
rect 3446 4358 3447 4364
rect 3451 4358 3452 4364
rect 3446 4354 3452 4358
rect 3446 4350 3447 4354
rect 3451 4350 3452 4354
rect 3446 4346 3452 4350
rect 3446 4342 3447 4346
rect 3451 4342 3452 4346
rect 3446 4338 3452 4342
rect 3446 4334 3447 4338
rect 3451 4334 3452 4338
rect 3446 4330 3452 4334
rect 3446 4326 3447 4330
rect 3451 4326 3452 4330
rect 3446 4322 3452 4326
rect 3446 4318 3447 4322
rect 3451 4318 3452 4322
rect 3446 4314 3452 4318
rect 3446 4310 3447 4314
rect 3451 4310 3452 4314
rect 3446 4306 3452 4310
rect 3446 4302 3447 4306
rect 3451 4302 3452 4306
rect 3446 4298 3452 4302
rect 3446 4294 3447 4298
rect 3451 4294 3452 4298
rect 3446 4290 3452 4294
rect 3446 4286 3447 4290
rect 3451 4286 3452 4290
rect 3446 4282 3452 4286
rect 3446 4278 3447 4282
rect 3451 4278 3452 4282
rect 3446 4274 3452 4278
rect 3446 4270 3447 4274
rect 3451 4270 3452 4274
rect 3446 4266 3452 4270
rect 3446 4262 3447 4266
rect 3451 4262 3452 4266
rect 3446 4258 3452 4262
rect 3446 4254 3447 4258
rect 3451 4254 3452 4258
rect 3446 4250 3452 4254
rect 3446 4246 3447 4250
rect 3451 4246 3452 4250
rect 3446 4245 3452 4246
<< pdcontact >>
rect 3393 4290 3397 4364
rect 3393 4246 3397 4268
rect 3405 4358 3409 4364
rect 3405 4350 3409 4354
rect 3405 4342 3409 4346
rect 3405 4334 3409 4338
rect 3405 4326 3409 4330
rect 3405 4318 3409 4322
rect 3405 4310 3409 4314
rect 3405 4302 3409 4306
rect 3405 4294 3409 4298
rect 3405 4286 3409 4290
rect 3405 4278 3409 4282
rect 3405 4270 3409 4274
rect 3405 4262 3409 4266
rect 3405 4254 3409 4258
rect 3405 4246 3409 4250
rect 3414 4246 3418 4364
rect 3426 4358 3430 4364
rect 3426 4350 3430 4354
rect 3426 4342 3430 4346
rect 3426 4334 3430 4338
rect 3426 4326 3430 4330
rect 3426 4318 3430 4322
rect 3426 4310 3430 4314
rect 3426 4302 3430 4306
rect 3426 4294 3430 4298
rect 3426 4286 3430 4290
rect 3426 4278 3430 4282
rect 3426 4270 3430 4274
rect 3426 4262 3430 4266
rect 3426 4254 3430 4258
rect 3426 4246 3430 4250
rect 3435 4246 3439 4364
rect 3447 4358 3451 4364
rect 3447 4350 3451 4354
rect 3447 4342 3451 4346
rect 3447 4334 3451 4338
rect 3447 4326 3451 4330
rect 3447 4318 3451 4322
rect 3447 4310 3451 4314
rect 3447 4302 3451 4306
rect 3447 4294 3451 4298
rect 3447 4286 3451 4290
rect 3447 4278 3451 4282
rect 3447 4270 3451 4274
rect 3447 4262 3451 4266
rect 3447 4254 3451 4258
rect 3447 4246 3451 4250
<< nsubstratencontact >>
rect 3463 4250 3508 4358
<< polysilicon >>
rect 3215 4369 3221 4374
rect 3398 4372 3446 4373
rect 3398 4367 3399 4372
rect 3445 4367 3446 4372
rect 3398 4366 3446 4367
rect 3398 4365 3404 4366
rect 3419 4365 3425 4366
rect 3440 4365 3446 4366
rect 3808 4358 3814 4363
rect 3398 4244 3404 4245
rect 3419 4244 3425 4245
rect 3440 4244 3446 4245
rect 3398 4243 3446 4244
rect 3398 4238 3399 4243
rect 3430 4238 3446 4243
rect 3398 4237 3446 4238
<< polycontact >>
rect 3399 4367 3445 4372
rect 3399 4238 3430 4243
<< metal1 >>
rect 1182 4528 1244 4529
rect 1013 4390 1053 4496
rect 1070 4404 1086 4496
rect 1159 4487 1244 4528
rect 1175 4486 1244 4487
rect 1198 4452 1244 4486
rect 1544 4474 1560 4507
rect 2018 4482 2034 4504
rect 1250 4404 1560 4474
rect 2006 4473 2047 4482
rect 1070 4393 1096 4404
rect 1244 4400 1560 4404
rect 1244 4393 1737 4397
rect 1013 4272 1101 4390
rect 1252 4381 1737 4393
rect 1289 4316 1737 4381
rect 1576 3948 1737 4316
rect 1981 4056 2072 4473
rect 2865 4067 2904 4500
rect 2910 4383 2948 4502
rect 3182 4463 3200 4464
rect 3182 4462 3346 4463
rect 3440 4462 3456 4511
rect 3182 4447 3456 4462
rect 3857 4460 3897 4489
rect 2910 4357 3176 4383
rect 3182 4364 3200 4447
rect 3344 4446 3456 4447
rect 3782 4418 3793 4419
rect 3782 4388 3784 4418
rect 3791 4388 3793 4418
rect 3414 4364 3418 4367
rect 2910 4343 3121 4357
rect 2910 4330 3058 4343
rect 3451 4358 3507 4359
rect 3451 4250 3463 4358
rect 3782 4354 3793 4388
rect 3817 4382 3897 4460
rect 3817 4346 3853 4382
rect 2865 4064 3051 4067
rect 1979 4007 2838 4056
rect 2865 4034 3214 4064
rect 3236 4007 3289 4246
rect 3414 4243 3418 4246
rect 3355 4240 3399 4243
rect 3355 4226 3356 4240
rect 3370 4238 3399 4240
rect 3435 4242 3439 4246
rect 3370 4226 3424 4238
rect 3435 4234 3458 4242
rect 3914 4238 3930 4505
rect 3355 4225 3424 4226
rect 3431 4097 3458 4234
rect 3826 4236 3930 4238
rect 3826 4206 3897 4236
rect 3927 4206 3930 4236
rect 3826 4202 3930 4206
rect 3431 4095 3635 4097
rect 3431 4061 3638 4095
rect 3991 4090 4031 4494
rect 4049 4404 4135 4405
rect 4045 4388 4492 4404
rect 4045 4366 4467 4388
rect 3431 4060 3635 4061
rect 3771 4051 4031 4090
rect 1979 3962 3289 4007
rect 2769 3961 3289 3962
rect 1576 3947 3599 3948
rect 4049 3947 4134 4366
rect 1576 3847 4134 3947
rect 4209 3991 4491 4031
rect 1409 3831 3376 3832
rect 1409 3817 3360 3831
rect 3375 3817 3376 3831
rect 4209 3830 4265 3991
rect 1409 3816 3376 3817
rect 1409 2034 1425 3816
rect 510 2018 1425 2034
rect 1437 3788 3587 3794
rect 1437 3721 3546 3788
rect 3578 3721 3587 3788
rect 3973 3780 4265 3830
rect 4374 3914 4491 3930
rect 1437 3716 3587 3721
rect 510 1558 528 1560
rect 504 1549 528 1558
rect 509 1544 528 1549
rect 573 1473 585 1485
rect 502 1443 585 1473
rect 1437 606 1515 3716
rect 3889 3682 3925 3684
rect 3889 3681 3930 3682
rect 1561 3679 3930 3681
rect 1561 3585 3898 3679
rect 1561 3584 3925 3585
rect 1561 1075 1658 3584
rect 3889 3583 3925 3584
rect 3974 3527 4024 3780
rect 4374 3756 4452 3914
rect 4086 3663 4452 3756
rect 4089 3335 4158 3663
rect 4309 3440 4491 3456
rect 4013 3293 4158 3335
rect 4310 3212 4349 3440
rect 4014 3176 4349 3212
rect 4013 3054 4279 3089
rect 3699 3031 3770 3043
rect 3699 2871 3743 3031
rect 3752 2960 4215 3027
rect 4249 2982 4279 3054
rect 4249 2966 4491 2982
rect 3983 2959 4215 2960
rect 4158 2949 4215 2959
rect 4158 2909 4491 2949
rect 3699 2869 4311 2871
rect 3699 2864 4312 2869
rect 3700 2808 4312 2864
rect 4229 2526 4312 2808
rect 4229 2508 4483 2526
rect 4229 2492 4491 2508
rect 4229 2471 4483 2492
rect 4457 2034 4484 2037
rect 4457 2018 4490 2034
rect 4457 2017 4484 2018
rect 4447 1961 4490 2001
rect 1561 1064 1564 1075
rect 1655 1064 1658 1075
rect 1561 1061 1658 1064
rect 1070 547 1521 606
rect 1070 508 1086 547
rect 1544 531 1554 1056
rect 4388 596 4490 612
rect 1544 512 1557 531
rect 1574 524 1661 535
rect 1621 510 1661 524
rect 4388 510 4404 596
<< m2contact >>
rect 3784 4388 3791 4418
rect 3216 4368 3220 4372
rect 3393 4268 3397 4290
rect 3405 4354 3409 4358
rect 3405 4346 3409 4350
rect 3405 4338 3409 4342
rect 3405 4330 3409 4334
rect 3405 4322 3409 4326
rect 3405 4314 3409 4318
rect 3405 4306 3409 4310
rect 3405 4298 3409 4302
rect 3405 4290 3409 4294
rect 3405 4282 3409 4286
rect 3405 4274 3409 4278
rect 3405 4266 3409 4270
rect 3405 4258 3409 4262
rect 3405 4250 3409 4254
rect 3426 4354 3430 4358
rect 3426 4346 3430 4350
rect 3426 4338 3430 4342
rect 3426 4330 3430 4334
rect 3426 4322 3430 4326
rect 3426 4314 3430 4318
rect 3426 4306 3430 4310
rect 3426 4298 3430 4302
rect 3426 4290 3430 4294
rect 3426 4282 3430 4286
rect 3426 4274 3430 4278
rect 3426 4266 3430 4270
rect 3426 4258 3430 4262
rect 3426 4250 3430 4254
rect 3447 4354 3451 4358
rect 3447 4346 3451 4350
rect 3447 4338 3451 4342
rect 3447 4330 3451 4334
rect 3447 4322 3451 4326
rect 3447 4314 3451 4318
rect 3447 4306 3451 4310
rect 3447 4298 3451 4302
rect 3447 4290 3451 4294
rect 3447 4282 3451 4286
rect 3447 4274 3451 4278
rect 3447 4266 3451 4270
rect 3447 4258 3451 4262
rect 3447 4250 3451 4254
rect 3809 4358 3813 4362
rect 3040 4095 3044 4099
rect 3356 4226 3370 4240
rect 3897 4206 3927 4236
rect 3360 3817 3375 3831
rect 3546 3721 3578 3788
rect 3898 3585 3926 3679
rect 1564 1064 1655 1075
rect 1562 525 1569 561
<< metal2 >>
rect 3485 4491 3513 4492
rect 2492 4476 2508 4491
rect 2452 3560 2543 4476
rect 2966 4417 2982 4491
rect 2966 4400 3228 4417
rect 2966 4399 3037 4400
rect 3212 4372 3227 4400
rect 3212 4368 3216 4372
rect 3220 4368 3227 4372
rect 3212 4364 3227 4368
rect 3473 4364 3513 4491
rect 4388 4477 4404 4487
rect 3405 4358 3513 4364
rect 3409 4354 3426 4358
rect 3430 4354 3447 4358
rect 3451 4354 3513 4358
rect 3405 4350 3513 4354
rect 3409 4346 3426 4350
rect 3430 4346 3447 4350
rect 3451 4346 3513 4350
rect 3405 4342 3513 4346
rect 3409 4338 3426 4342
rect 3430 4338 3447 4342
rect 3451 4338 3513 4342
rect 3405 4334 3513 4338
rect 3409 4330 3426 4334
rect 3430 4330 3447 4334
rect 3451 4330 3513 4334
rect 3405 4326 3513 4330
rect 3409 4322 3426 4326
rect 3430 4322 3447 4326
rect 3451 4322 3513 4326
rect 3405 4318 3513 4322
rect 3409 4314 3426 4318
rect 3430 4314 3447 4318
rect 3451 4314 3513 4318
rect 3405 4310 3513 4314
rect 3409 4306 3426 4310
rect 3430 4306 3447 4310
rect 3451 4306 3513 4310
rect 3405 4302 3513 4306
rect 3409 4298 3426 4302
rect 3430 4298 3447 4302
rect 3451 4298 3513 4302
rect 3405 4294 3513 4298
rect 3106 4290 3395 4291
rect 3409 4290 3426 4294
rect 3430 4290 3447 4294
rect 3451 4290 3513 4294
rect 3106 4268 3393 4290
rect 3405 4286 3513 4290
rect 3409 4282 3426 4286
rect 3430 4282 3447 4286
rect 3451 4282 3513 4286
rect 3405 4278 3513 4282
rect 3409 4274 3426 4278
rect 3430 4274 3447 4278
rect 3451 4274 3513 4278
rect 3405 4270 3513 4274
rect 3106 4267 3395 4268
rect 3106 4266 3149 4267
rect 3409 4266 3426 4270
rect 3430 4266 3447 4270
rect 3451 4266 3513 4270
rect 3106 4172 3126 4266
rect 3405 4262 3513 4266
rect 3409 4258 3426 4262
rect 3430 4258 3447 4262
rect 3451 4258 3513 4262
rect 3405 4254 3513 4258
rect 3409 4250 3426 4254
rect 3430 4250 3447 4254
rect 3451 4250 3513 4254
rect 3405 4246 3513 4250
rect 3534 4419 3599 4420
rect 3534 4418 3793 4419
rect 3534 4388 3784 4418
rect 3791 4388 3793 4418
rect 3534 4387 3793 4388
rect 3039 4159 3126 4172
rect 3355 4240 3371 4241
rect 3355 4226 3356 4240
rect 3370 4226 3371 4240
rect 3039 4099 3056 4159
rect 3039 4095 3040 4099
rect 3044 4095 3056 4099
rect 3039 4092 3056 4095
rect 3355 3831 3371 4226
rect 3355 3817 3360 3831
rect 3355 3816 3371 3817
rect 3534 3788 3599 4387
rect 3805 4366 4404 4477
rect 3805 4362 3816 4366
rect 3805 4358 3809 4362
rect 3813 4358 3816 4362
rect 3805 4354 3816 4358
rect 3898 4236 3930 4246
rect 3927 4206 3930 4236
rect 3534 3721 3546 3788
rect 3578 3721 3599 3788
rect 3534 3714 3599 3721
rect 3898 3876 3930 4206
rect 3898 3679 3931 3876
rect 3926 3586 3931 3679
rect 2452 3513 3738 3560
rect 2452 3478 3782 3513
rect 2452 3477 3738 3478
rect 2452 3476 2543 3477
rect 925 2467 2513 2468
rect 866 2401 2513 2467
rect 866 636 924 2401
rect 523 613 924 636
rect 509 599 924 613
rect 1561 1075 1658 1080
rect 1561 1064 1564 1075
rect 1655 1064 1658 1075
rect 509 597 923 599
rect 523 585 923 597
rect 1561 561 1658 1064
rect 569 529 612 543
rect 596 510 611 529
rect 1561 525 1562 561
rect 1569 525 1658 561
rect 1561 524 1658 525
use blankpad  blankpad_11
timestamp 1259953556
transform -1 0 841 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_0
timestamp 1259953556
transform -1 0 1315 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_1
timestamp 1259953556
transform -1 0 1789 0 -1 5000
box -2 0 476 513
use inpad  inpad_9
timestamp 1259953556
transform -1 0 2263 0 -1 5000
box -2 0 476 513
use inpad  inpad_8
timestamp 1259953556
transform -1 0 2737 0 -1 5000
box -2 0 476 513
use inpad  inpad_7
timestamp 1259953556
transform -1 0 3211 0 -1 5000
box -2 0 476 513
use inpad  inpad_6
timestamp 1259953556
transform -1 0 3685 0 -1 5000
box -2 0 476 513
use inpad  inpad_5
timestamp 1259953556
transform -1 0 4159 0 -1 5000
box -2 0 476 513
use inpadp2  inpadp2_0
timestamp 1418813110
transform -1 0 4633 0 -1 5000
box -2 0 476 513
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 4487
box 0 0 5000 513
use blankpad  blankpad_27
timestamp 1259953556
transform 0 1 0 -1 0 4633
box -2 0 476 513
use inpad  inpad_12
timestamp 1259953556
transform 0 1 0 -1 0 4159
box -2 0 476 513
use inpad  inpad_13
timestamp 1259953556
transform 0 1 0 -1 0 3685
box -2 0 476 513
use inpad  inpad_14
timestamp 1259953556
transform 0 1 0 -1 0 3211
box -2 0 476 513
use inpad  inpad_15
timestamp 1259953556
transform 0 1 0 -1 0 2737
box -2 0 476 513
use inpad  inpad_16
timestamp 1259953556
transform 0 1 0 -1 0 2263
box -2 0 476 513
use 2-OR  2-OR_0
timestamp 1418434502
transform -1 0 1392 0 -1 4250
box 147 -223 302 -14
use Opamp  Opamp_0
timestamp 1418826157
transform 1 0 3221 0 1 4072
box -193 -11 77 303
use Opamp  Opamp_1
timestamp 1418826157
transform 1 0 3814 0 1 4062
box -193 -11 77 303
use DAC  DAC_0
timestamp 1418788810
transform -1 0 4009 0 -1 3535
box -14 4 257 511
use inpad  inpad_3
timestamp 1259953556
transform 0 -1 5000 1 0 4159
box -2 0 476 513
use inpad  inpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 3685
box -2 0 476 513
use inpad  inpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 3211
box -2 0 476 513
use inpad  inpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 2737
box -2 0 476 513
use inpad  inpad_11
timestamp 1259953556
transform 0 -1 5000 1 0 2263
box -2 0 476 513
use 50K_resistor  50K_resistor_0
timestamp 1418811347
transform -1 0 4601 0 -1 2225
box 143 188 207 270
use 50K_resistor  50K_resistor_1
timestamp 1418811347
transform -1 0 727 0 -1 1746
box 143 188 207 270
use inpad  inpad_17
timestamp 1259953556
transform 0 1 0 -1 0 1789
box -2 0 476 513
use inpad  inpad_18
timestamp 1259953556
transform 0 1 0 -1 0 1315
box -2 0 476 513
use Inductor  Inductor_0
timestamp 1418825699
transform 1 0 572 0 1 537
box -1 -1 3800 3800
use inpad  inpad_19
timestamp 1259953556
transform 0 -1 5000 1 0 1789
box -2 0 476 513
use blankpad  blankpad_8
timestamp 1259953556
transform 0 -1 5000 1 0 1315
box -2 0 476 513
use blankpad  blankpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 841
box -2 0 476 513
use 2_200K_resistors  2_200K_resistors_0
timestamp 1418810336
transform 0 -1 1838 1 0 354
box 170 181 703 290
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 367
box 2 2 513 4264
use barepad  barepad_3
timestamp 1259953556
transform 0 1 0 -1 0 841
box -2 0 476 513
use barepad  barepad_2
timestamp 1259953556
transform 1 0 367 0 1 0
box -2 0 476 513
use inpad  inpad_10
timestamp 1259953556
transform 1 0 841 0 1 0
box -2 0 476 513
use inpad  inpad_4
timestamp 1259953556
transform 1 0 1315 0 1 0
box -2 0 476 513
use blankpad  blankpad_25
timestamp 1259953556
transform 1 0 1789 0 1 0
box -2 0 476 513
use blankpad  blankpad_24
timestamp 1259953556
transform 1 0 2263 0 1 0
box -2 0 476 513
use blankpad  blankpad_23
timestamp 1259953556
transform 1 0 2737 0 1 0
box -2 0 476 513
use blankpad  blankpad_22
timestamp 1259953556
transform 1 0 3211 0 1 0
box -2 0 476 513
use blankpad  blankpad_21
timestamp 1259953556
transform 1 0 3685 0 1 0
box -2 0 476 513
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 4487 0 1 367
box 0 2 511 4264
use barepad  barepad_0
timestamp 1259953556
transform 0 -1 5000 1 0 367
box -2 0 476 513
use barepad  barepad_1
timestamp 1259953556
transform 1 0 4159 0 1 0
box -2 0 476 513
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 5000 513
<< end >>
