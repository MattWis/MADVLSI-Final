magic
tech scmos
timestamp 1418434502
<< nwell >>
rect 147 -150 302 -14
<< ntransistor >>
rect 162 -162 164 -156
rect 172 -162 174 -156
rect 180 -162 182 -156
rect 197 -216 199 -156
rect 214 -216 216 -156
rect 222 -216 224 -156
rect 230 -216 232 -156
rect 238 -216 240 -156
rect 246 -216 248 -156
rect 254 -216 256 -156
rect 262 -216 264 -156
rect 270 -216 272 -156
rect 278 -216 280 -156
rect 286 -216 288 -156
<< ptransistor >>
rect 163 -141 165 -135
rect 168 -141 170 -135
rect 178 -144 180 -132
rect 197 -141 199 -21
rect 216 -141 218 -21
rect 224 -141 226 -21
rect 232 -141 234 -21
rect 240 -141 242 -21
rect 248 -141 250 -21
rect 256 -141 258 -21
rect 264 -141 266 -21
rect 272 -141 274 -21
rect 280 -141 282 -21
rect 288 -141 290 -21
<< ndiffusion >>
rect 156 -157 162 -156
rect 156 -161 157 -157
rect 161 -161 162 -157
rect 156 -162 162 -161
rect 164 -157 172 -156
rect 164 -161 165 -157
rect 171 -161 172 -157
rect 164 -162 172 -161
rect 174 -157 180 -156
rect 174 -161 175 -157
rect 179 -161 180 -157
rect 174 -162 180 -161
rect 182 -157 188 -156
rect 182 -161 183 -157
rect 187 -161 188 -157
rect 182 -162 188 -161
rect 191 -157 197 -156
rect 191 -161 192 -157
rect 196 -161 197 -157
rect 165 -166 171 -162
rect 191 -165 197 -161
rect 191 -169 192 -165
rect 196 -169 197 -165
rect 191 -173 197 -169
rect 191 -177 192 -173
rect 196 -177 197 -173
rect 191 -181 197 -177
rect 191 -191 192 -181
rect 196 -191 197 -181
rect 191 -195 197 -191
rect 191 -199 192 -195
rect 196 -199 197 -195
rect 191 -203 197 -199
rect 191 -207 192 -203
rect 196 -207 197 -203
rect 191 -211 197 -207
rect 191 -215 192 -211
rect 196 -215 197 -211
rect 191 -216 197 -215
rect 199 -157 205 -156
rect 199 -215 200 -157
rect 204 -215 205 -157
rect 199 -216 205 -215
rect 208 -157 214 -156
rect 208 -161 209 -157
rect 213 -161 214 -157
rect 208 -165 214 -161
rect 208 -169 209 -165
rect 213 -169 214 -165
rect 208 -173 214 -169
rect 208 -177 209 -173
rect 213 -177 214 -173
rect 208 -181 214 -177
rect 208 -191 209 -181
rect 213 -191 214 -181
rect 208 -195 214 -191
rect 208 -199 209 -195
rect 213 -199 214 -195
rect 208 -203 214 -199
rect 208 -207 209 -203
rect 213 -207 214 -203
rect 208 -211 214 -207
rect 208 -215 209 -211
rect 213 -215 214 -211
rect 208 -216 214 -215
rect 216 -157 222 -156
rect 216 -215 217 -157
rect 221 -215 222 -157
rect 216 -216 222 -215
rect 224 -157 230 -156
rect 224 -161 225 -157
rect 229 -161 230 -157
rect 224 -165 230 -161
rect 224 -169 225 -165
rect 229 -169 230 -165
rect 224 -173 230 -169
rect 224 -177 225 -173
rect 229 -177 230 -173
rect 224 -181 230 -177
rect 224 -191 225 -181
rect 229 -191 230 -181
rect 224 -195 230 -191
rect 224 -199 225 -195
rect 229 -199 230 -195
rect 224 -203 230 -199
rect 224 -207 225 -203
rect 229 -207 230 -203
rect 224 -211 230 -207
rect 224 -215 225 -211
rect 229 -215 230 -211
rect 224 -216 230 -215
rect 232 -157 238 -156
rect 232 -215 233 -157
rect 237 -215 238 -157
rect 232 -216 238 -215
rect 240 -157 246 -156
rect 240 -161 241 -157
rect 245 -161 246 -157
rect 240 -165 246 -161
rect 240 -169 241 -165
rect 245 -169 246 -165
rect 240 -173 246 -169
rect 240 -177 241 -173
rect 245 -177 246 -173
rect 240 -181 246 -177
rect 240 -191 241 -181
rect 245 -191 246 -181
rect 240 -195 246 -191
rect 240 -199 241 -195
rect 245 -199 246 -195
rect 240 -203 246 -199
rect 240 -207 241 -203
rect 245 -207 246 -203
rect 240 -211 246 -207
rect 240 -215 241 -211
rect 245 -215 246 -211
rect 240 -216 246 -215
rect 248 -157 254 -156
rect 248 -215 249 -157
rect 253 -215 254 -157
rect 248 -216 254 -215
rect 256 -157 262 -156
rect 256 -161 257 -157
rect 261 -161 262 -157
rect 256 -165 262 -161
rect 256 -169 257 -165
rect 261 -169 262 -165
rect 256 -173 262 -169
rect 256 -177 257 -173
rect 261 -177 262 -173
rect 256 -181 262 -177
rect 256 -191 257 -181
rect 261 -191 262 -181
rect 256 -195 262 -191
rect 256 -199 257 -195
rect 261 -199 262 -195
rect 256 -203 262 -199
rect 256 -207 257 -203
rect 261 -207 262 -203
rect 256 -211 262 -207
rect 256 -215 257 -211
rect 261 -215 262 -211
rect 256 -216 262 -215
rect 264 -157 270 -156
rect 264 -215 265 -157
rect 269 -215 270 -157
rect 264 -216 270 -215
rect 272 -157 278 -156
rect 272 -161 273 -157
rect 277 -161 278 -157
rect 272 -165 278 -161
rect 272 -169 273 -165
rect 277 -169 278 -165
rect 272 -173 278 -169
rect 272 -177 273 -173
rect 277 -177 278 -173
rect 272 -181 278 -177
rect 272 -191 273 -181
rect 277 -191 278 -181
rect 272 -195 278 -191
rect 272 -199 273 -195
rect 277 -199 278 -195
rect 272 -203 278 -199
rect 272 -207 273 -203
rect 277 -207 278 -203
rect 272 -211 278 -207
rect 272 -215 273 -211
rect 277 -215 278 -211
rect 272 -216 278 -215
rect 280 -157 286 -156
rect 280 -215 281 -157
rect 285 -215 286 -157
rect 280 -216 286 -215
rect 288 -157 294 -156
rect 288 -161 289 -157
rect 293 -161 294 -157
rect 288 -165 294 -161
rect 288 -169 289 -165
rect 293 -169 294 -165
rect 288 -173 294 -169
rect 288 -177 289 -173
rect 293 -177 294 -173
rect 288 -181 294 -177
rect 288 -191 289 -181
rect 293 -191 294 -181
rect 288 -195 294 -191
rect 288 -199 289 -195
rect 293 -199 294 -195
rect 288 -203 294 -199
rect 288 -207 289 -203
rect 293 -207 294 -203
rect 288 -211 294 -207
rect 288 -215 289 -211
rect 293 -215 294 -211
rect 288 -216 294 -215
<< pdiffusion >>
rect 191 -24 197 -21
rect 191 -28 192 -24
rect 196 -28 197 -24
rect 191 -32 197 -28
rect 191 -36 192 -32
rect 196 -36 197 -32
rect 191 -40 197 -36
rect 191 -44 192 -40
rect 196 -44 197 -40
rect 191 -48 197 -44
rect 191 -52 192 -48
rect 196 -52 197 -48
rect 191 -56 197 -52
rect 191 -60 192 -56
rect 196 -60 197 -56
rect 191 -64 197 -60
rect 191 -68 192 -64
rect 196 -68 197 -64
rect 191 -72 197 -68
rect 191 -76 192 -72
rect 196 -76 197 -72
rect 191 -80 197 -76
rect 191 -84 192 -80
rect 196 -84 197 -80
rect 191 -88 197 -84
rect 191 -92 192 -88
rect 196 -92 197 -88
rect 191 -96 197 -92
rect 191 -100 192 -96
rect 196 -100 197 -96
rect 191 -104 197 -100
rect 191 -108 192 -104
rect 196 -108 197 -104
rect 191 -112 197 -108
rect 191 -116 192 -112
rect 196 -116 197 -112
rect 191 -120 197 -116
rect 191 -124 192 -120
rect 196 -124 197 -120
rect 191 -128 197 -124
rect 191 -132 192 -128
rect 196 -132 197 -128
rect 175 -135 178 -132
rect 153 -136 163 -135
rect 153 -140 158 -136
rect 162 -140 163 -136
rect 153 -141 163 -140
rect 165 -141 168 -135
rect 170 -136 178 -135
rect 170 -140 172 -136
rect 176 -140 178 -136
rect 170 -141 178 -140
rect 175 -144 178 -141
rect 180 -136 186 -132
rect 180 -140 181 -136
rect 185 -140 186 -136
rect 180 -144 186 -140
rect 191 -136 197 -132
rect 191 -140 192 -136
rect 196 -140 197 -136
rect 191 -141 197 -140
rect 199 -22 205 -21
rect 199 -140 200 -22
rect 204 -140 205 -22
rect 199 -141 205 -140
rect 210 -22 216 -21
rect 210 -28 211 -22
rect 215 -28 216 -22
rect 210 -32 216 -28
rect 210 -36 211 -32
rect 215 -36 216 -32
rect 210 -40 216 -36
rect 210 -44 211 -40
rect 215 -44 216 -40
rect 210 -48 216 -44
rect 210 -52 211 -48
rect 215 -52 216 -48
rect 210 -56 216 -52
rect 210 -60 211 -56
rect 215 -60 216 -56
rect 210 -64 216 -60
rect 210 -68 211 -64
rect 215 -68 216 -64
rect 210 -72 216 -68
rect 210 -76 211 -72
rect 215 -76 216 -72
rect 210 -80 216 -76
rect 210 -84 211 -80
rect 215 -84 216 -80
rect 210 -88 216 -84
rect 210 -92 211 -88
rect 215 -92 216 -88
rect 210 -96 216 -92
rect 210 -100 211 -96
rect 215 -100 216 -96
rect 210 -104 216 -100
rect 210 -108 211 -104
rect 215 -108 216 -104
rect 210 -112 216 -108
rect 210 -116 211 -112
rect 215 -116 216 -112
rect 210 -120 216 -116
rect 210 -124 211 -120
rect 215 -124 216 -120
rect 210 -128 216 -124
rect 210 -132 211 -128
rect 215 -132 216 -128
rect 210 -136 216 -132
rect 210 -140 211 -136
rect 215 -140 216 -136
rect 210 -141 216 -140
rect 218 -22 224 -21
rect 218 -140 219 -22
rect 223 -140 224 -22
rect 218 -141 224 -140
rect 226 -22 232 -21
rect 226 -28 227 -22
rect 231 -28 232 -22
rect 226 -32 232 -28
rect 226 -36 227 -32
rect 231 -36 232 -32
rect 226 -40 232 -36
rect 226 -44 227 -40
rect 231 -44 232 -40
rect 226 -48 232 -44
rect 226 -52 227 -48
rect 231 -52 232 -48
rect 226 -56 232 -52
rect 226 -60 227 -56
rect 231 -60 232 -56
rect 226 -64 232 -60
rect 226 -68 227 -64
rect 231 -68 232 -64
rect 226 -72 232 -68
rect 226 -76 227 -72
rect 231 -76 232 -72
rect 226 -80 232 -76
rect 226 -84 227 -80
rect 231 -84 232 -80
rect 226 -88 232 -84
rect 226 -92 227 -88
rect 231 -92 232 -88
rect 226 -96 232 -92
rect 226 -100 227 -96
rect 231 -100 232 -96
rect 226 -104 232 -100
rect 226 -108 227 -104
rect 231 -108 232 -104
rect 226 -112 232 -108
rect 226 -116 227 -112
rect 231 -116 232 -112
rect 226 -120 232 -116
rect 226 -124 227 -120
rect 231 -124 232 -120
rect 226 -128 232 -124
rect 226 -132 227 -128
rect 231 -132 232 -128
rect 226 -136 232 -132
rect 226 -140 227 -136
rect 231 -140 232 -136
rect 226 -141 232 -140
rect 234 -22 240 -21
rect 234 -140 235 -22
rect 239 -140 240 -22
rect 234 -141 240 -140
rect 242 -22 248 -21
rect 242 -28 243 -22
rect 247 -28 248 -22
rect 242 -32 248 -28
rect 242 -36 243 -32
rect 247 -36 248 -32
rect 242 -40 248 -36
rect 242 -44 243 -40
rect 247 -44 248 -40
rect 242 -48 248 -44
rect 242 -52 243 -48
rect 247 -52 248 -48
rect 242 -56 248 -52
rect 242 -60 243 -56
rect 247 -60 248 -56
rect 242 -64 248 -60
rect 242 -68 243 -64
rect 247 -68 248 -64
rect 242 -72 248 -68
rect 242 -76 243 -72
rect 247 -76 248 -72
rect 242 -80 248 -76
rect 242 -84 243 -80
rect 247 -84 248 -80
rect 242 -88 248 -84
rect 242 -92 243 -88
rect 247 -92 248 -88
rect 242 -96 248 -92
rect 242 -100 243 -96
rect 247 -100 248 -96
rect 242 -104 248 -100
rect 242 -108 243 -104
rect 247 -108 248 -104
rect 242 -112 248 -108
rect 242 -116 243 -112
rect 247 -116 248 -112
rect 242 -120 248 -116
rect 242 -124 243 -120
rect 247 -124 248 -120
rect 242 -128 248 -124
rect 242 -132 243 -128
rect 247 -132 248 -128
rect 242 -136 248 -132
rect 242 -140 243 -136
rect 247 -140 248 -136
rect 242 -141 248 -140
rect 250 -22 256 -21
rect 250 -140 251 -22
rect 255 -140 256 -22
rect 250 -141 256 -140
rect 258 -22 264 -21
rect 258 -28 259 -22
rect 263 -28 264 -22
rect 258 -32 264 -28
rect 258 -36 259 -32
rect 263 -36 264 -32
rect 258 -40 264 -36
rect 258 -44 259 -40
rect 263 -44 264 -40
rect 258 -48 264 -44
rect 258 -52 259 -48
rect 263 -52 264 -48
rect 258 -56 264 -52
rect 258 -60 259 -56
rect 263 -60 264 -56
rect 258 -64 264 -60
rect 258 -68 259 -64
rect 263 -68 264 -64
rect 258 -72 264 -68
rect 258 -76 259 -72
rect 263 -76 264 -72
rect 258 -80 264 -76
rect 258 -84 259 -80
rect 263 -84 264 -80
rect 258 -88 264 -84
rect 258 -92 259 -88
rect 263 -92 264 -88
rect 258 -96 264 -92
rect 258 -100 259 -96
rect 263 -100 264 -96
rect 258 -104 264 -100
rect 258 -108 259 -104
rect 263 -108 264 -104
rect 258 -112 264 -108
rect 258 -116 259 -112
rect 263 -116 264 -112
rect 258 -120 264 -116
rect 258 -124 259 -120
rect 263 -124 264 -120
rect 258 -128 264 -124
rect 258 -132 259 -128
rect 263 -132 264 -128
rect 258 -136 264 -132
rect 258 -140 259 -136
rect 263 -140 264 -136
rect 258 -141 264 -140
rect 266 -22 272 -21
rect 266 -140 267 -22
rect 271 -140 272 -22
rect 266 -141 272 -140
rect 274 -22 280 -21
rect 274 -28 275 -22
rect 279 -28 280 -22
rect 274 -32 280 -28
rect 274 -36 275 -32
rect 279 -36 280 -32
rect 274 -40 280 -36
rect 274 -44 275 -40
rect 279 -44 280 -40
rect 274 -48 280 -44
rect 274 -52 275 -48
rect 279 -52 280 -48
rect 274 -56 280 -52
rect 274 -60 275 -56
rect 279 -60 280 -56
rect 274 -64 280 -60
rect 274 -68 275 -64
rect 279 -68 280 -64
rect 274 -72 280 -68
rect 274 -76 275 -72
rect 279 -76 280 -72
rect 274 -80 280 -76
rect 274 -84 275 -80
rect 279 -84 280 -80
rect 274 -88 280 -84
rect 274 -92 275 -88
rect 279 -92 280 -88
rect 274 -96 280 -92
rect 274 -100 275 -96
rect 279 -100 280 -96
rect 274 -104 280 -100
rect 274 -108 275 -104
rect 279 -108 280 -104
rect 274 -112 280 -108
rect 274 -116 275 -112
rect 279 -116 280 -112
rect 274 -120 280 -116
rect 274 -124 275 -120
rect 279 -124 280 -120
rect 274 -128 280 -124
rect 274 -132 275 -128
rect 279 -132 280 -128
rect 274 -136 280 -132
rect 274 -140 275 -136
rect 279 -140 280 -136
rect 274 -141 280 -140
rect 282 -22 288 -21
rect 282 -140 283 -22
rect 287 -140 288 -22
rect 282 -141 288 -140
rect 290 -22 296 -21
rect 290 -28 291 -22
rect 295 -28 296 -22
rect 290 -32 296 -28
rect 290 -36 291 -32
rect 295 -36 296 -32
rect 290 -40 296 -36
rect 290 -44 291 -40
rect 295 -44 296 -40
rect 290 -48 296 -44
rect 290 -52 291 -48
rect 295 -52 296 -48
rect 290 -56 296 -52
rect 290 -60 291 -56
rect 295 -60 296 -56
rect 290 -64 296 -60
rect 290 -68 291 -64
rect 295 -68 296 -64
rect 290 -72 296 -68
rect 290 -76 291 -72
rect 295 -76 296 -72
rect 290 -80 296 -76
rect 290 -84 291 -80
rect 295 -84 296 -80
rect 290 -88 296 -84
rect 290 -92 291 -88
rect 295 -92 296 -88
rect 290 -96 296 -92
rect 290 -100 291 -96
rect 295 -100 296 -96
rect 290 -104 296 -100
rect 290 -108 291 -104
rect 295 -108 296 -104
rect 290 -112 296 -108
rect 290 -116 291 -112
rect 295 -116 296 -112
rect 290 -120 296 -116
rect 290 -124 291 -120
rect 295 -124 296 -120
rect 290 -128 296 -124
rect 290 -132 291 -128
rect 295 -132 296 -128
rect 290 -136 296 -132
rect 290 -140 291 -136
rect 295 -140 296 -136
rect 290 -141 296 -140
<< ndcontact >>
rect 157 -161 161 -157
rect 165 -161 171 -157
rect 175 -161 179 -157
rect 183 -161 187 -157
rect 192 -161 196 -157
rect 192 -169 196 -165
rect 192 -177 196 -173
rect 192 -191 196 -181
rect 192 -199 196 -195
rect 192 -207 196 -203
rect 192 -215 196 -211
rect 200 -215 204 -157
rect 209 -161 213 -157
rect 209 -169 213 -165
rect 209 -177 213 -173
rect 209 -191 213 -181
rect 209 -199 213 -195
rect 209 -207 213 -203
rect 209 -215 213 -211
rect 217 -215 221 -157
rect 225 -161 229 -157
rect 225 -169 229 -165
rect 225 -177 229 -173
rect 225 -191 229 -181
rect 225 -199 229 -195
rect 225 -207 229 -203
rect 225 -215 229 -211
rect 233 -215 237 -157
rect 241 -161 245 -157
rect 241 -169 245 -165
rect 241 -177 245 -173
rect 241 -191 245 -181
rect 241 -199 245 -195
rect 241 -207 245 -203
rect 241 -215 245 -211
rect 249 -215 253 -157
rect 257 -161 261 -157
rect 257 -169 261 -165
rect 257 -177 261 -173
rect 257 -191 261 -181
rect 257 -199 261 -195
rect 257 -207 261 -203
rect 257 -215 261 -211
rect 265 -215 269 -157
rect 273 -161 277 -157
rect 273 -169 277 -165
rect 273 -177 277 -173
rect 273 -191 277 -181
rect 273 -199 277 -195
rect 273 -207 277 -203
rect 273 -215 277 -211
rect 281 -215 285 -157
rect 289 -161 293 -157
rect 289 -169 293 -165
rect 289 -177 293 -173
rect 289 -191 293 -181
rect 289 -199 293 -195
rect 289 -207 293 -203
rect 289 -215 293 -211
<< pdcontact >>
rect 192 -28 196 -24
rect 192 -36 196 -32
rect 192 -44 196 -40
rect 192 -52 196 -48
rect 192 -60 196 -56
rect 192 -68 196 -64
rect 192 -76 196 -72
rect 192 -84 196 -80
rect 192 -92 196 -88
rect 192 -100 196 -96
rect 192 -108 196 -104
rect 192 -116 196 -112
rect 192 -124 196 -120
rect 192 -132 196 -128
rect 158 -140 162 -136
rect 172 -140 176 -136
rect 181 -140 185 -136
rect 192 -140 196 -136
rect 200 -140 204 -22
rect 211 -28 215 -22
rect 211 -36 215 -32
rect 211 -44 215 -40
rect 211 -52 215 -48
rect 211 -60 215 -56
rect 211 -68 215 -64
rect 211 -76 215 -72
rect 211 -84 215 -80
rect 211 -92 215 -88
rect 211 -100 215 -96
rect 211 -108 215 -104
rect 211 -116 215 -112
rect 211 -124 215 -120
rect 211 -132 215 -128
rect 211 -140 215 -136
rect 219 -140 223 -22
rect 227 -28 231 -22
rect 227 -36 231 -32
rect 227 -44 231 -40
rect 227 -52 231 -48
rect 227 -60 231 -56
rect 227 -68 231 -64
rect 227 -76 231 -72
rect 227 -84 231 -80
rect 227 -92 231 -88
rect 227 -100 231 -96
rect 227 -108 231 -104
rect 227 -116 231 -112
rect 227 -124 231 -120
rect 227 -132 231 -128
rect 227 -140 231 -136
rect 235 -140 239 -22
rect 243 -28 247 -22
rect 243 -36 247 -32
rect 243 -44 247 -40
rect 243 -52 247 -48
rect 243 -60 247 -56
rect 243 -68 247 -64
rect 243 -76 247 -72
rect 243 -84 247 -80
rect 243 -92 247 -88
rect 243 -100 247 -96
rect 243 -108 247 -104
rect 243 -116 247 -112
rect 243 -124 247 -120
rect 243 -132 247 -128
rect 243 -140 247 -136
rect 251 -140 255 -22
rect 259 -28 263 -22
rect 259 -36 263 -32
rect 259 -44 263 -40
rect 259 -52 263 -48
rect 259 -60 263 -56
rect 259 -68 263 -64
rect 259 -76 263 -72
rect 259 -84 263 -80
rect 259 -92 263 -88
rect 259 -100 263 -96
rect 259 -108 263 -104
rect 259 -116 263 -112
rect 259 -124 263 -120
rect 259 -132 263 -128
rect 259 -140 263 -136
rect 267 -140 271 -22
rect 275 -28 279 -22
rect 275 -36 279 -32
rect 275 -44 279 -40
rect 275 -52 279 -48
rect 275 -60 279 -56
rect 275 -68 279 -64
rect 275 -76 279 -72
rect 275 -84 279 -80
rect 275 -92 279 -88
rect 275 -100 279 -96
rect 275 -108 279 -104
rect 275 -116 279 -112
rect 275 -124 279 -120
rect 275 -132 279 -128
rect 275 -140 279 -136
rect 283 -140 287 -22
rect 291 -28 295 -22
rect 291 -36 295 -32
rect 291 -44 295 -40
rect 291 -52 295 -48
rect 291 -60 295 -56
rect 291 -68 295 -64
rect 291 -76 295 -72
rect 291 -84 295 -80
rect 291 -92 295 -88
rect 291 -100 295 -96
rect 291 -108 295 -104
rect 291 -116 295 -112
rect 291 -124 295 -120
rect 291 -132 295 -128
rect 291 -140 295 -136
<< psubstratepcontact >>
rect 148 -216 191 -170
<< nsubstratencontact >>
rect 150 -128 191 -22
<< polysilicon >>
rect 216 -15 290 -14
rect 216 -19 217 -15
rect 289 -19 290 -15
rect 197 -21 199 -19
rect 216 -20 290 -19
rect 216 -21 218 -20
rect 224 -21 226 -20
rect 232 -21 234 -20
rect 240 -21 242 -20
rect 248 -21 250 -20
rect 256 -21 258 -20
rect 264 -21 266 -20
rect 272 -21 274 -20
rect 280 -21 282 -20
rect 288 -21 290 -20
rect 178 -132 180 -130
rect 163 -135 165 -133
rect 168 -135 170 -133
rect 163 -149 165 -141
rect 168 -142 170 -141
rect 168 -143 174 -142
rect 168 -147 169 -143
rect 173 -147 174 -143
rect 197 -142 199 -141
rect 216 -142 218 -141
rect 224 -142 226 -141
rect 232 -142 234 -141
rect 240 -142 242 -141
rect 248 -142 250 -141
rect 256 -142 258 -141
rect 264 -142 266 -141
rect 272 -142 274 -141
rect 280 -142 282 -141
rect 288 -142 290 -141
rect 168 -148 174 -147
rect 158 -150 165 -149
rect 158 -154 159 -150
rect 163 -154 165 -150
rect 158 -155 165 -154
rect 171 -155 174 -148
rect 178 -149 180 -144
rect 193 -147 199 -142
rect 177 -150 183 -149
rect 177 -154 178 -150
rect 182 -154 183 -150
rect 177 -155 183 -154
rect 193 -151 194 -147
rect 198 -151 199 -147
rect 193 -155 199 -151
rect 210 -143 294 -142
rect 210 -154 211 -143
rect 215 -154 294 -143
rect 210 -155 294 -154
rect 162 -156 164 -155
rect 172 -156 174 -155
rect 180 -156 182 -155
rect 197 -156 199 -155
rect 214 -156 216 -155
rect 222 -156 224 -155
rect 230 -156 232 -155
rect 238 -156 240 -155
rect 246 -156 248 -155
rect 254 -156 256 -155
rect 262 -156 264 -155
rect 270 -156 272 -155
rect 278 -156 280 -155
rect 286 -156 288 -155
rect 162 -164 164 -162
rect 172 -164 174 -162
rect 180 -164 182 -162
rect 197 -218 199 -216
rect 214 -217 216 -216
rect 222 -217 224 -216
rect 230 -217 232 -216
rect 238 -217 240 -216
rect 246 -217 248 -216
rect 254 -217 256 -216
rect 262 -217 264 -216
rect 270 -217 272 -216
rect 278 -217 280 -216
rect 286 -217 288 -216
rect 214 -218 288 -217
rect 214 -222 215 -218
rect 287 -222 288 -218
rect 214 -223 288 -222
<< polycontact >>
rect 217 -19 289 -15
rect 169 -147 173 -143
rect 159 -154 163 -150
rect 178 -154 182 -150
rect 194 -151 198 -147
rect 211 -154 215 -143
rect 215 -222 287 -218
<< metal1 >>
rect 147 -22 192 -21
rect 147 -128 150 -22
rect 191 -128 192 -22
rect 147 -133 192 -128
rect 170 -136 178 -133
rect 170 -140 172 -136
rect 176 -140 178 -136
rect 147 -147 169 -143
rect 185 -147 189 -136
rect 204 -140 205 -22
rect 210 -140 211 -22
rect 223 -140 224 -22
rect 239 -140 240 -22
rect 255 -140 256 -22
rect 271 -140 272 -22
rect 287 -140 288 -22
rect 200 -143 205 -140
rect 219 -142 224 -140
rect 218 -143 224 -142
rect 235 -143 240 -140
rect 251 -143 256 -140
rect 267 -143 272 -140
rect 283 -143 288 -140
rect 200 -144 211 -143
rect 147 -154 159 -150
rect 166 -154 178 -150
rect 185 -151 194 -147
rect 166 -157 170 -154
rect 185 -157 189 -151
rect 201 -154 211 -144
rect 218 -154 300 -143
rect 200 -157 205 -154
rect 218 -157 222 -154
rect 234 -157 238 -154
rect 250 -157 254 -154
rect 266 -157 270 -154
rect 282 -157 286 -154
rect 147 -161 157 -157
rect 187 -161 189 -157
rect 147 -169 161 -161
rect 175 -169 179 -161
rect 147 -170 192 -169
rect 147 -216 148 -170
rect 191 -215 192 -170
rect 204 -215 205 -157
rect 221 -215 222 -157
rect 237 -215 238 -157
rect 253 -215 254 -157
rect 269 -215 270 -157
rect 285 -215 286 -157
rect 191 -216 196 -215
rect 147 -217 196 -216
<< m2contact >>
rect 192 -32 196 -28
rect 192 -40 196 -36
rect 192 -48 196 -44
rect 192 -56 196 -52
rect 192 -64 196 -60
rect 192 -72 196 -68
rect 192 -80 196 -76
rect 192 -88 196 -84
rect 192 -96 196 -92
rect 192 -104 196 -100
rect 192 -112 196 -108
rect 192 -120 196 -116
rect 192 -128 196 -124
rect 192 -136 196 -132
rect 154 -140 158 -136
rect 211 -32 215 -28
rect 211 -40 215 -36
rect 211 -48 215 -44
rect 211 -56 215 -52
rect 211 -64 215 -60
rect 211 -72 215 -68
rect 211 -80 215 -76
rect 211 -88 215 -84
rect 211 -96 215 -92
rect 211 -104 215 -100
rect 211 -112 215 -108
rect 211 -120 215 -116
rect 211 -128 215 -124
rect 211 -136 215 -132
rect 227 -32 231 -28
rect 227 -40 231 -36
rect 227 -48 231 -44
rect 227 -56 231 -52
rect 227 -64 231 -60
rect 227 -72 231 -68
rect 227 -80 231 -76
rect 227 -88 231 -84
rect 227 -96 231 -92
rect 227 -104 231 -100
rect 227 -112 231 -108
rect 227 -120 231 -116
rect 227 -128 231 -124
rect 227 -136 231 -132
rect 243 -32 247 -28
rect 243 -40 247 -36
rect 243 -48 247 -44
rect 243 -56 247 -52
rect 243 -64 247 -60
rect 243 -72 247 -68
rect 243 -80 247 -76
rect 243 -88 247 -84
rect 243 -96 247 -92
rect 243 -104 247 -100
rect 243 -112 247 -108
rect 243 -120 247 -116
rect 243 -128 247 -124
rect 243 -136 247 -132
rect 259 -32 263 -28
rect 259 -40 263 -36
rect 259 -48 263 -44
rect 259 -56 263 -52
rect 259 -64 263 -60
rect 259 -72 263 -68
rect 259 -80 263 -76
rect 259 -88 263 -84
rect 259 -96 263 -92
rect 259 -104 263 -100
rect 259 -112 263 -108
rect 259 -120 263 -116
rect 259 -128 263 -124
rect 259 -136 263 -132
rect 275 -32 279 -28
rect 275 -40 279 -36
rect 275 -48 279 -44
rect 275 -56 279 -52
rect 275 -64 279 -60
rect 275 -72 279 -68
rect 275 -80 279 -76
rect 275 -88 279 -84
rect 275 -96 279 -92
rect 275 -104 279 -100
rect 275 -112 279 -108
rect 275 -120 279 -116
rect 275 -128 279 -124
rect 275 -136 279 -132
rect 291 -32 295 -28
rect 291 -40 295 -36
rect 291 -48 295 -44
rect 291 -56 295 -52
rect 291 -64 295 -60
rect 291 -72 295 -68
rect 291 -80 295 -76
rect 291 -88 295 -84
rect 291 -96 295 -92
rect 291 -104 295 -100
rect 291 -112 295 -108
rect 291 -120 295 -116
rect 291 -128 295 -124
rect 291 -136 295 -132
rect 166 -165 170 -161
rect 192 -165 196 -161
rect 192 -173 196 -169
rect 192 -181 196 -177
rect 192 -195 196 -191
rect 192 -203 196 -199
rect 192 -211 196 -207
rect 209 -165 213 -161
rect 209 -173 213 -169
rect 209 -181 213 -177
rect 209 -195 213 -191
rect 209 -203 213 -199
rect 209 -211 213 -207
rect 225 -165 229 -161
rect 225 -173 229 -169
rect 225 -181 229 -177
rect 225 -195 229 -191
rect 225 -203 229 -199
rect 225 -211 229 -207
rect 241 -165 245 -161
rect 241 -173 245 -169
rect 241 -181 245 -177
rect 241 -195 245 -191
rect 241 -203 245 -199
rect 241 -211 245 -207
rect 257 -165 261 -161
rect 257 -173 261 -169
rect 257 -181 261 -177
rect 257 -195 261 -191
rect 257 -203 261 -199
rect 257 -211 261 -207
rect 273 -165 277 -161
rect 273 -173 277 -169
rect 273 -181 277 -177
rect 273 -195 277 -191
rect 273 -203 277 -199
rect 273 -211 277 -207
rect 289 -165 293 -161
rect 289 -173 293 -169
rect 289 -181 293 -177
rect 289 -195 293 -191
rect 289 -203 293 -199
rect 289 -211 293 -207
<< metal2 >>
rect 192 -28 302 -22
rect 196 -32 211 -28
rect 215 -32 227 -28
rect 231 -32 243 -28
rect 247 -32 259 -28
rect 263 -32 275 -28
rect 279 -32 291 -28
rect 295 -32 302 -28
rect 192 -36 302 -32
rect 196 -40 211 -36
rect 215 -40 227 -36
rect 231 -40 243 -36
rect 247 -40 259 -36
rect 263 -40 275 -36
rect 279 -40 291 -36
rect 295 -40 302 -36
rect 192 -44 302 -40
rect 196 -48 211 -44
rect 215 -48 227 -44
rect 231 -48 243 -44
rect 247 -48 259 -44
rect 263 -48 275 -44
rect 279 -48 291 -44
rect 295 -48 302 -44
rect 192 -52 302 -48
rect 196 -56 211 -52
rect 215 -56 227 -52
rect 231 -56 243 -52
rect 247 -56 259 -52
rect 263 -56 275 -52
rect 279 -56 291 -52
rect 295 -56 302 -52
rect 192 -60 302 -56
rect 196 -64 211 -60
rect 215 -64 227 -60
rect 231 -64 243 -60
rect 247 -64 259 -60
rect 263 -64 275 -60
rect 279 -64 291 -60
rect 295 -64 302 -60
rect 192 -68 302 -64
rect 196 -72 211 -68
rect 215 -72 227 -68
rect 231 -72 243 -68
rect 247 -72 259 -68
rect 263 -72 275 -68
rect 279 -72 291 -68
rect 295 -72 302 -68
rect 192 -76 302 -72
rect 196 -80 211 -76
rect 215 -80 227 -76
rect 231 -80 243 -76
rect 247 -80 259 -76
rect 263 -80 275 -76
rect 279 -80 291 -76
rect 295 -80 302 -76
rect 192 -84 302 -80
rect 196 -88 211 -84
rect 215 -88 227 -84
rect 231 -88 243 -84
rect 247 -88 259 -84
rect 263 -88 275 -84
rect 279 -88 291 -84
rect 295 -88 302 -84
rect 192 -92 302 -88
rect 196 -96 211 -92
rect 215 -96 227 -92
rect 231 -96 243 -92
rect 247 -96 259 -92
rect 263 -96 275 -92
rect 279 -96 291 -92
rect 295 -96 302 -92
rect 192 -100 302 -96
rect 196 -104 211 -100
rect 215 -104 227 -100
rect 231 -104 243 -100
rect 247 -104 259 -100
rect 263 -104 275 -100
rect 279 -104 291 -100
rect 295 -104 302 -100
rect 192 -108 302 -104
rect 196 -112 211 -108
rect 215 -112 227 -108
rect 231 -112 243 -108
rect 247 -112 259 -108
rect 263 -112 275 -108
rect 279 -112 291 -108
rect 295 -112 302 -108
rect 192 -116 302 -112
rect 196 -120 211 -116
rect 215 -120 227 -116
rect 231 -120 243 -116
rect 247 -120 259 -116
rect 263 -120 275 -116
rect 279 -120 291 -116
rect 295 -120 302 -116
rect 192 -124 302 -120
rect 196 -128 211 -124
rect 215 -128 227 -124
rect 231 -128 243 -124
rect 247 -128 259 -124
rect 263 -128 275 -124
rect 279 -128 291 -124
rect 295 -128 302 -124
rect 192 -132 302 -128
rect 196 -136 211 -132
rect 215 -136 227 -132
rect 231 -136 243 -132
rect 247 -136 259 -132
rect 263 -136 275 -132
rect 279 -136 291 -132
rect 295 -136 302 -132
rect 158 -147 162 -136
rect 192 -140 302 -136
rect 158 -151 170 -147
rect 166 -157 170 -151
rect 165 -161 170 -157
rect 192 -161 293 -157
rect 196 -165 209 -161
rect 213 -165 225 -161
rect 229 -165 241 -161
rect 245 -165 257 -161
rect 261 -165 273 -161
rect 277 -165 289 -161
rect 192 -169 293 -165
rect 196 -173 209 -169
rect 213 -173 225 -169
rect 229 -173 241 -169
rect 245 -173 257 -169
rect 261 -173 273 -169
rect 277 -173 289 -169
rect 192 -177 293 -173
rect 196 -181 209 -177
rect 213 -181 225 -177
rect 229 -181 241 -177
rect 245 -181 257 -177
rect 261 -181 273 -177
rect 277 -181 289 -177
rect 192 -191 293 -181
rect 196 -195 209 -191
rect 213 -195 225 -191
rect 229 -195 241 -191
rect 245 -195 257 -191
rect 261 -195 273 -191
rect 277 -195 289 -191
rect 192 -199 293 -195
rect 196 -203 209 -199
rect 213 -203 225 -199
rect 229 -203 241 -199
rect 245 -203 257 -199
rect 261 -203 273 -199
rect 277 -203 289 -199
rect 192 -207 293 -203
rect 196 -211 209 -207
rect 213 -211 225 -207
rect 229 -211 241 -207
rect 245 -211 257 -207
rect 261 -211 273 -207
rect 277 -211 289 -207
rect 192 -215 293 -211
<< labels >>
rlabel metal1 155 -154 159 -150 1 B
rlabel metal1 155 -147 169 -143 1 A
rlabel metal1 218 -154 300 -143 1 Z
rlabel metal1 154 -161 157 -157 1 Gnd
<< end >>
