magic
tech scmos
timestamp 1418788065
<< electrode >>
rect 159 486 164 488
rect 159 434 164 436
rect 159 425 164 427
rect 159 373 164 375
rect 159 364 164 366
rect 159 312 164 314
rect 159 303 164 305
rect 159 251 164 253
rect 159 242 164 244
rect 159 190 164 192
rect 159 181 164 183
rect 159 129 164 131
rect 159 120 164 122
rect 159 68 164 70
rect 159 55 164 57
rect 159 3 164 5
<< genericpoly2contact >>
rect 159 488 164 492
rect 159 427 164 434
rect 159 366 164 373
rect 159 305 164 312
rect 159 244 164 251
rect 159 183 164 190
rect 159 122 164 129
rect 159 57 164 68
rect 159 -1 164 3
<< metal1 >>
rect 155 497 177 500
rect 155 490 177 493
rect 158 489 177 490
rect 158 487 165 489
rect 158 432 165 435
rect 155 429 165 432
rect 158 426 165 429
rect 158 371 165 374
rect 155 368 165 371
rect 158 365 165 368
rect 158 310 165 313
rect 155 307 165 310
rect 158 304 165 307
rect 158 249 165 252
rect 155 246 165 249
rect 158 243 165 246
rect 158 188 165 191
rect 155 185 165 188
rect 158 182 165 185
rect 158 127 165 130
rect 155 124 165 127
rect 158 121 165 124
rect 158 66 165 69
rect 155 63 165 66
rect 158 56 165 63
rect 171 11 177 14
rect 158 -4 165 4
rect 155 -7 177 -4
<< m2contact >>
rect 167 11 171 15
<< metal2 >>
rect 155 11 167 15
<< high_resist >>
rect 157 436 159 486
rect 164 436 166 486
rect 157 375 159 425
rect 164 375 166 425
rect 157 314 159 364
rect 164 314 166 364
rect 157 253 159 303
rect 164 253 166 303
rect 157 192 159 242
rect 164 192 166 242
rect 157 131 159 181
rect 164 131 166 181
rect 157 70 159 120
rect 164 70 166 120
rect 157 5 159 55
rect 164 5 166 55
<< poly2_high_resist >>
rect 159 436 164 486
rect 159 375 164 425
rect 159 314 164 364
rect 159 253 164 303
rect 159 192 164 242
rect 159 131 164 181
rect 159 70 164 120
rect 159 5 164 55
<< labels >>
rlabel metal1 175 11 177 14 7 DAC_Output
rlabel metal1 175 -7 177 -4 8 gnd
rlabel metal1 175 497 177 500 6 vdd
rlabel metal1 175 489 177 493 7 Rin
rlabel metal1 155 429 156 432 3 bit6
rlabel metal1 155 368 156 371 3 bit5
rlabel metal1 155 307 156 310 3 bit4
rlabel metal1 155 246 156 249 3 bit3
rlabel metal1 155 185 156 188 3 bit2
rlabel metal1 155 124 156 127 3 bit1
rlabel metal1 155 63 156 66 3 bit0
rlabel metal1 155 490 156 493 3 bit7
<< end >>
