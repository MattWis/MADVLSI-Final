magic
tech scmos
timestamp 1415734409
<< nwell >>
rect 69 -109 207 42
rect 97 -117 134 -109
<< ntransistor >>
rect 187 -128 193 -122
rect 86 -249 92 -129
rect 98 -249 104 -129
rect 122 -249 128 -129
rect 146 -249 152 -129
rect 158 -249 164 -129
rect 170 -249 176 -129
<< ptransistor >>
rect 86 -101 92 19
rect 98 -101 104 19
rect 140 -101 146 19
rect 152 -101 158 19
rect 176 -101 182 19
rect 113 -108 119 -102
<< ndiffusion >>
rect 187 -117 193 -116
rect 187 -121 188 -117
rect 192 -121 193 -117
rect 187 -122 193 -121
rect 187 -129 193 -128
rect 80 -232 86 -129
rect 80 -236 81 -232
rect 85 -236 86 -232
rect 80 -249 86 -236
rect 92 -243 98 -129
rect 92 -247 93 -243
rect 97 -247 98 -243
rect 92 -249 98 -247
rect 104 -133 110 -129
rect 104 -137 105 -133
rect 109 -137 110 -133
rect 104 -249 110 -137
rect 116 -134 122 -129
rect 116 -138 117 -134
rect 121 -138 122 -134
rect 116 -249 122 -138
rect 128 -232 134 -129
rect 128 -236 129 -232
rect 133 -236 134 -232
rect 128 -249 134 -236
rect 140 -133 146 -129
rect 140 -137 141 -133
rect 145 -137 146 -133
rect 140 -249 146 -137
rect 152 -232 158 -129
rect 152 -236 153 -232
rect 157 -236 158 -232
rect 152 -249 158 -236
rect 164 -243 170 -129
rect 164 -247 165 -243
rect 169 -247 170 -243
rect 164 -249 170 -247
rect 176 -131 182 -129
rect 176 -135 177 -131
rect 181 -135 182 -131
rect 176 -249 182 -135
rect 187 -133 188 -129
rect 192 -133 193 -129
rect 187 -138 193 -133
<< pdiffusion >>
rect 80 -94 86 19
rect 80 -98 81 -94
rect 85 -98 86 -94
rect 80 -101 86 -98
rect 92 17 98 19
rect 92 13 93 17
rect 97 13 98 17
rect 92 -101 98 13
rect 104 -75 110 19
rect 104 -79 105 -75
rect 109 -79 110 -75
rect 104 -101 110 -79
rect 134 -32 140 19
rect 134 -36 135 -32
rect 139 -36 140 -32
rect 113 -97 119 -92
rect 113 -101 114 -97
rect 118 -101 119 -97
rect 134 -101 140 -36
rect 146 3 152 19
rect 146 -1 147 3
rect 151 -1 152 3
rect 146 -101 152 -1
rect 158 17 164 19
rect 158 13 159 17
rect 163 13 164 17
rect 158 -101 164 13
rect 170 3 176 19
rect 170 -1 171 3
rect 175 -1 176 3
rect 170 -101 176 -1
rect 182 17 188 19
rect 182 13 183 17
rect 187 13 188 17
rect 182 -94 188 13
rect 182 -98 183 -94
rect 187 -98 188 -94
rect 182 -101 188 -98
rect 113 -102 119 -101
rect 113 -109 119 -108
rect 113 -113 114 -109
rect 118 -113 119 -109
rect 113 -114 119 -113
<< ndcontact >>
rect 188 -121 192 -117
rect 81 -236 85 -232
rect 93 -247 97 -243
rect 105 -137 109 -133
rect 117 -138 121 -134
rect 129 -236 133 -232
rect 141 -137 145 -133
rect 153 -236 157 -232
rect 165 -247 169 -243
rect 177 -135 181 -131
rect 188 -133 192 -129
<< pdcontact >>
rect 81 -98 85 -94
rect 93 13 97 17
rect 105 -79 109 -75
rect 135 -36 139 -32
rect 114 -101 118 -97
rect 147 -1 151 3
rect 159 13 163 17
rect 171 -1 175 3
rect 183 13 187 17
rect 183 -98 187 -94
rect 114 -113 118 -109
<< psubstratepcontact >>
rect 188 -142 192 -138
rect 78 -265 82 -261
<< nsubstratencontact >>
rect 114 -92 118 -88
<< polysilicon >>
rect 152 25 182 26
rect 86 20 104 22
rect 152 21 177 25
rect 181 21 182 25
rect 86 19 92 20
rect 98 19 104 20
rect 140 19 146 21
rect 152 20 182 21
rect 152 19 158 20
rect 176 19 182 20
rect 86 -102 92 -101
rect 98 -102 104 -101
rect 140 -102 146 -101
rect 86 -103 113 -102
rect 86 -107 87 -103
rect 91 -107 113 -103
rect 86 -108 113 -107
rect 119 -108 125 -102
rect 140 -106 141 -102
rect 145 -106 146 -102
rect 152 -103 158 -101
rect 176 -103 182 -101
rect 140 -107 146 -106
rect 122 -121 164 -117
rect 122 -124 128 -121
rect 86 -128 104 -126
rect 86 -129 92 -128
rect 98 -129 104 -128
rect 122 -128 123 -124
rect 127 -128 128 -124
rect 122 -129 128 -128
rect 146 -124 152 -123
rect 146 -128 147 -124
rect 151 -128 152 -124
rect 146 -129 152 -128
rect 158 -129 164 -121
rect 170 -128 187 -122
rect 193 -128 195 -122
rect 170 -129 176 -128
rect 86 -250 92 -249
rect 98 -250 104 -249
rect 86 -251 104 -250
rect 122 -251 128 -249
rect 146 -251 152 -249
rect 158 -251 164 -249
rect 86 -255 87 -251
rect 91 -254 104 -251
rect 170 -254 176 -249
rect 91 -255 176 -254
rect 86 -256 176 -255
rect 99 -260 176 -256
<< polycontact >>
rect 177 21 181 25
rect 87 -107 91 -103
rect 141 -106 145 -102
rect 123 -128 127 -124
rect 147 -128 151 -124
rect 87 -255 91 -251
<< metal1 >>
rect 158 34 194 35
rect 158 29 207 34
rect 158 18 164 29
rect 192 28 207 29
rect 176 25 188 26
rect 176 21 177 25
rect 181 21 188 25
rect 176 20 188 21
rect 69 17 164 18
rect 69 12 93 17
rect 97 13 159 17
rect 163 13 164 17
rect 97 12 164 13
rect 182 17 188 20
rect 182 13 183 17
rect 187 13 207 17
rect 182 12 207 13
rect 146 3 176 4
rect 146 -1 147 3
rect 151 -1 171 3
rect 175 -1 176 3
rect 146 -2 176 -1
rect 134 -36 135 -31
rect 139 -36 146 -31
rect 134 -37 146 -36
rect 104 -75 128 -74
rect 104 -79 105 -75
rect 109 -79 128 -75
rect 104 -80 128 -79
rect 113 -88 119 -87
rect 113 -92 114 -88
rect 118 -92 119 -88
rect 113 -93 119 -92
rect 80 -94 92 -93
rect 80 -98 81 -94
rect 85 -98 92 -94
rect 80 -99 92 -98
rect 86 -103 92 -99
rect 113 -101 114 -93
rect 118 -101 119 -93
rect 113 -102 119 -101
rect 86 -107 87 -103
rect 91 -107 92 -103
rect 86 -132 92 -107
rect 113 -109 119 -108
rect 113 -113 114 -109
rect 118 -113 119 -109
rect 113 -123 119 -113
rect 122 -114 128 -80
rect 140 -101 146 -37
rect 182 -94 193 -93
rect 182 -98 183 -94
rect 187 -98 193 -94
rect 182 -99 193 -98
rect 140 -102 170 -101
rect 140 -106 141 -102
rect 145 -106 170 -102
rect 140 -107 170 -106
rect 122 -120 138 -114
rect 132 -123 138 -120
rect 113 -124 128 -123
rect 113 -128 123 -124
rect 127 -128 128 -124
rect 113 -129 128 -128
rect 132 -124 152 -123
rect 132 -128 147 -124
rect 151 -128 152 -124
rect 132 -129 152 -128
rect 86 -133 110 -132
rect 86 -137 105 -133
rect 109 -137 110 -133
rect 86 -138 110 -137
rect 116 -134 122 -129
rect 116 -138 117 -134
rect 121 -138 122 -134
rect 116 -197 122 -138
rect 140 -133 146 -129
rect 140 -137 141 -133
rect 145 -137 146 -133
rect 164 -130 170 -107
rect 187 -117 193 -99
rect 187 -121 188 -117
rect 192 -121 193 -117
rect 187 -122 193 -121
rect 164 -131 182 -130
rect 164 -135 177 -131
rect 181 -135 182 -131
rect 164 -136 182 -135
rect 140 -187 146 -137
rect 187 -137 188 -129
rect 192 -137 193 -129
rect 187 -138 193 -137
rect 187 -142 188 -138
rect 192 -142 193 -138
rect 187 -143 193 -142
rect 140 -193 207 -187
rect 116 -203 207 -197
rect 196 -214 207 -208
rect 80 -232 86 -231
rect 80 -236 81 -232
rect 85 -236 86 -232
rect 80 -250 86 -236
rect 128 -232 158 -231
rect 128 -236 129 -232
rect 133 -236 153 -232
rect 157 -236 158 -232
rect 128 -237 158 -236
rect 93 -243 165 -241
rect 196 -241 202 -214
rect 97 -247 165 -243
rect 169 -247 202 -241
rect 69 -251 92 -250
rect 69 -255 87 -251
rect 91 -255 92 -251
rect 69 -256 92 -255
rect 100 -260 106 -247
rect 69 -261 106 -260
rect 69 -265 78 -261
rect 82 -265 106 -261
rect 69 -266 106 -265
<< m2contact >>
rect 93 9 97 13
rect 135 -32 139 -28
rect 114 -97 118 -93
rect 188 -137 192 -133
rect 165 -243 169 -239
<< metal2 >>
rect 92 13 119 14
rect 92 9 93 13
rect 97 9 119 13
rect 92 8 119 9
rect 113 -93 119 8
rect 134 -1 207 5
rect 134 -28 140 -1
rect 134 -32 135 -28
rect 139 -32 140 -28
rect 134 -37 140 -32
rect 113 -97 114 -93
rect 118 -97 119 -93
rect 113 -98 119 -97
rect 187 -133 193 -132
rect 187 -137 188 -133
rect 192 -137 193 -133
rect 187 -238 193 -137
rect 164 -239 193 -238
rect 164 -243 165 -239
rect 169 -243 193 -239
rect 164 -244 193 -243
<< labels >>
rlabel metal1 192 28 207 34 1 Vdd
rlabel metal1 187 12 207 17 1 Vbp
rlabel metal2 134 -1 207 5 1 Vcp
rlabel metal1 140 -193 207 -187 1 Vcn
rlabel metal1 116 -203 207 -197 1 Vbn
rlabel metal1 69 -256 87 -250 1 Iin
rlabel metal1 69 12 93 18 1 Vdd
rlabel metal1 86 -138 92 -107 1 Iip
<< end >>
