magic
tech scmos
timestamp 1418333373
<< error_s >>
rect -317 282 -316 288
<< polysilicon >>
rect -363 295 -324 296
rect -363 291 -362 295
rect -325 291 -324 295
rect -363 290 -324 291
rect -363 289 -357 290
rect -351 289 -345 290
rect -330 289 -324 290
rect -363 168 -357 169
rect -351 168 -345 169
rect -330 168 -324 169
rect -363 167 -324 168
rect -363 163 -362 167
rect -347 163 -337 167
rect -325 163 -324 167
rect -363 162 -324 163
<< ndiffusion >>
rect -155 12 -139 26
<< pdiffusion >>
rect -369 288 -363 289
rect -369 170 -368 288
rect -364 170 -363 288
rect -369 169 -363 170
rect -357 288 -351 289
rect -357 282 -356 288
rect -352 282 -351 288
rect -357 278 -351 282
rect -357 274 -356 278
rect -352 274 -351 278
rect -357 270 -351 274
rect -357 266 -356 270
rect -352 266 -351 270
rect -357 262 -351 266
rect -357 258 -356 262
rect -352 258 -351 262
rect -357 254 -351 258
rect -357 250 -356 254
rect -352 250 -351 254
rect -357 246 -351 250
rect -357 242 -356 246
rect -352 242 -351 246
rect -357 238 -351 242
rect -357 234 -356 238
rect -352 234 -351 238
rect -357 230 -351 234
rect -357 226 -356 230
rect -352 226 -351 230
rect -357 222 -351 226
rect -357 218 -356 222
rect -352 218 -351 222
rect -357 214 -351 218
rect -357 210 -356 214
rect -352 210 -351 214
rect -357 206 -351 210
rect -357 202 -356 206
rect -352 202 -351 206
rect -357 198 -351 202
rect -357 194 -356 198
rect -352 194 -351 198
rect -357 190 -351 194
rect -357 186 -356 190
rect -352 186 -351 190
rect -357 182 -351 186
rect -357 178 -356 182
rect -352 178 -351 182
rect -357 174 -351 178
rect -357 170 -356 174
rect -352 170 -351 174
rect -357 169 -351 170
rect -345 288 -339 289
rect -345 170 -344 288
rect -340 170 -339 288
rect -345 169 -339 170
rect -336 288 -330 289
rect -336 282 -335 288
rect -331 282 -330 288
rect -336 278 -330 282
rect -336 274 -335 278
rect -331 274 -330 278
rect -336 270 -330 274
rect -336 266 -335 270
rect -331 266 -330 270
rect -336 262 -330 266
rect -336 258 -335 262
rect -331 258 -330 262
rect -336 254 -330 258
rect -336 250 -335 254
rect -331 250 -330 254
rect -336 246 -330 250
rect -336 242 -335 246
rect -331 242 -330 246
rect -336 238 -330 242
rect -336 234 -335 238
rect -331 234 -330 238
rect -336 230 -330 234
rect -336 226 -335 230
rect -331 226 -330 230
rect -336 222 -330 226
rect -336 218 -335 222
rect -331 218 -330 222
rect -336 214 -330 218
rect -336 210 -335 214
rect -331 210 -330 214
rect -336 206 -330 210
rect -336 202 -335 206
rect -331 202 -330 206
rect -336 198 -330 202
rect -336 194 -335 198
rect -331 194 -330 198
rect -336 190 -330 194
rect -336 186 -335 190
rect -331 186 -330 190
rect -336 182 -330 186
rect -336 178 -335 182
rect -331 178 -330 182
rect -336 174 -330 178
rect -336 170 -335 174
rect -331 170 -330 174
rect -336 169 -330 170
rect -324 288 -318 289
rect -324 170 -323 288
rect -319 170 -318 288
rect -324 169 -318 170
<< metal1 >>
rect -368 291 -362 295
rect -368 288 -360 291
rect -364 170 -360 288
rect -319 170 -314 270
rect -368 167 -360 170
rect -368 163 -362 167
rect -344 160 -340 170
rect -347 -6 -337 160
rect -322 14 -314 170
rect -157 13 -154 25
rect -347 -16 -92 -6
rect -102 -147 -92 -16
rect -60 -135 -47 -107
rect -102 -172 -72 -147
rect -64 -157 -47 -135
rect -64 -161 74 -157
rect -60 -182 74 -161
<< metal2 >>
rect -336 288 -276 289
rect -383 282 -276 288
rect -383 278 -356 282
rect -352 278 -335 282
rect -331 278 -276 282
rect -383 274 -331 278
rect -383 270 -356 274
rect -352 270 -335 274
rect -383 266 -331 270
rect -383 262 -356 266
rect -352 262 -335 266
rect -383 258 -331 262
rect -383 254 -356 258
rect -352 254 -335 258
rect -383 250 -331 254
rect -383 246 -356 250
rect -352 246 -335 250
rect -383 242 -331 246
rect -383 238 -356 242
rect -352 238 -335 242
rect -383 234 -331 238
rect -383 230 -356 234
rect -352 230 -335 234
rect -383 226 -331 230
rect -383 222 -356 226
rect -352 222 -335 226
rect -331 222 -38 224
rect -383 218 -38 222
rect -383 214 -356 218
rect -352 214 -335 218
rect -331 214 -38 218
rect -383 210 -38 214
rect -383 206 -356 210
rect -352 206 -335 210
rect -331 206 -38 210
rect -383 202 -38 206
rect -383 198 -356 202
rect -352 198 -335 202
rect -331 198 -38 202
rect -383 194 -38 198
rect -383 190 -356 194
rect -352 190 -335 194
rect -331 190 -38 194
rect -383 186 -38 190
rect -383 182 -356 186
rect -352 182 -335 186
rect -331 184 -38 186
rect -383 178 -331 182
rect -383 174 -356 178
rect -352 174 -335 178
rect -383 170 -331 174
rect -77 92 -38 184
rect -140 13 -93 25
rect -107 -107 -93 13
rect -107 -111 -64 -107
rect -107 -115 -60 -111
rect -107 -119 -64 -115
rect -107 -123 -60 -119
rect -107 -127 -64 -123
rect -107 -131 -60 -127
rect -107 -135 -64 -131
<< ptransistor >>
rect -363 169 -357 289
rect -351 169 -345 289
rect -330 169 -324 289
<< polycontact >>
rect -362 291 -325 295
rect -362 163 -347 167
rect -337 163 -325 167
<< ndcontact >>
rect -64 -115 -60 -111
rect -64 -123 -60 -119
rect -64 -131 -60 -127
<< pdcontact >>
rect -368 170 -364 288
rect -356 282 -352 288
rect -356 274 -352 278
rect -356 266 -352 270
rect -356 258 -352 262
rect -356 250 -352 254
rect -356 242 -352 246
rect -356 234 -352 238
rect -356 226 -352 230
rect -356 218 -352 222
rect -356 210 -352 214
rect -356 202 -352 206
rect -356 194 -352 198
rect -356 186 -352 190
rect -356 178 -352 182
rect -356 170 -352 174
rect -344 170 -340 288
rect -335 282 -331 288
rect -335 274 -331 278
rect -335 266 -331 270
rect -335 258 -331 262
rect -335 250 -331 254
rect -335 242 -331 246
rect -335 234 -331 238
rect -335 226 -331 230
rect -335 218 -331 222
rect -335 210 -331 214
rect -335 202 -331 206
rect -335 194 -331 198
rect -335 186 -331 190
rect -335 178 -331 182
rect -335 170 -331 174
rect -323 170 -319 288
<< m2contact >>
rect -356 278 -352 282
rect -356 270 -352 274
rect -356 262 -352 266
rect -356 254 -352 258
rect -356 246 -352 250
rect -356 238 -352 242
rect -356 230 -352 234
rect -356 222 -352 226
rect -356 214 -352 218
rect -356 206 -352 210
rect -356 198 -352 202
rect -356 190 -352 194
rect -356 182 -352 186
rect -356 174 -352 178
rect -335 278 -331 282
rect -335 270 -331 274
rect -335 262 -331 266
rect -335 254 -331 258
rect -335 246 -331 250
rect -335 238 -331 242
rect -335 230 -331 234
rect -335 222 -331 226
rect -335 214 -331 218
rect -335 206 -331 210
rect -335 198 -331 202
rect -335 190 -331 194
rect -335 182 -331 186
rect -335 174 -331 178
rect -154 13 -140 25
rect -64 -111 -60 -107
rect -64 -119 -60 -115
rect -64 -127 -60 -123
rect -64 -135 -60 -131
use Opamp  Opamp_0
timestamp 1418331768
transform 1 0 -124 0 1 15
box -193 -11 77 303
use Opamp  Opamp_1
timestamp 1418331768
transform 1 0 105 0 1 -171
box -193 -11 77 303
<< end >>
