magic
tech scmos
timestamp 1418333453
<< metal1 >>
rect -66 14 -9 47
rect -160 -11 -66 14
<< psubstratepcontact >>
rect -66 -11 -9 14
use Bias  Bias_0
timestamp 1415734409
transform 1 0 -262 0 1 255
box 69 -266 207 42
use FCDAmp  FCDAmp_0
timestamp 1414784736
transform 1 0 -28 0 1 92
box -27 -68 105 211
<< labels >>
rlabel metal1 -52 10 -37 47 1 Gnd
<< end >>
