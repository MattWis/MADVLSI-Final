magic
tech scmos
timestamp 1418814466
<< error_p >>
rect 1562 3681 1564 3682
<< error_s >>
rect 796 4679 797 4683
rect 802 4679 803 4683
rect 808 4679 809 4683
rect 814 4679 815 4683
rect 820 4679 821 4683
rect 826 4679 827 4683
rect 858 4679 859 4683
rect 864 4679 865 4683
rect 870 4679 871 4683
rect 876 4679 877 4683
rect 882 4679 883 4683
rect 888 4679 889 4683
rect 1270 4679 1271 4683
rect 1276 4679 1277 4683
rect 1282 4679 1283 4683
rect 1288 4679 1289 4683
rect 1294 4679 1295 4683
rect 1300 4679 1301 4683
rect 1332 4679 1333 4683
rect 1338 4679 1339 4683
rect 1344 4679 1345 4683
rect 1350 4679 1351 4683
rect 1356 4679 1357 4683
rect 1362 4679 1363 4683
rect 1744 4679 1745 4683
rect 1750 4679 1751 4683
rect 1756 4679 1757 4683
rect 1762 4679 1763 4683
rect 1768 4679 1769 4683
rect 1774 4679 1775 4683
rect 796 4667 797 4671
rect 802 4667 803 4671
rect 808 4667 809 4671
rect 814 4667 815 4671
rect 820 4667 821 4671
rect 826 4667 827 4671
rect 858 4667 859 4671
rect 864 4667 865 4671
rect 870 4667 871 4671
rect 876 4667 877 4671
rect 882 4667 883 4671
rect 888 4667 889 4671
rect 1270 4667 1271 4671
rect 1276 4667 1277 4671
rect 1282 4667 1283 4671
rect 1288 4667 1289 4671
rect 1294 4667 1295 4671
rect 1300 4667 1301 4671
rect 1332 4667 1333 4671
rect 1338 4667 1339 4671
rect 1344 4667 1345 4671
rect 1350 4667 1351 4671
rect 1356 4667 1357 4671
rect 1362 4667 1363 4671
rect 1744 4667 1745 4671
rect 1750 4667 1751 4671
rect 1756 4667 1757 4671
rect 1762 4667 1763 4671
rect 1768 4667 1769 4671
rect 1774 4667 1775 4671
rect 796 4655 797 4659
rect 802 4655 803 4659
rect 808 4655 809 4659
rect 814 4655 815 4659
rect 820 4655 821 4659
rect 826 4655 827 4659
rect 858 4655 859 4659
rect 864 4655 865 4659
rect 870 4655 871 4659
rect 876 4655 877 4659
rect 882 4655 883 4659
rect 888 4655 889 4659
rect 1270 4655 1271 4659
rect 1276 4655 1277 4659
rect 1282 4655 1283 4659
rect 1288 4655 1289 4659
rect 1294 4655 1295 4659
rect 1300 4655 1301 4659
rect 1332 4655 1333 4659
rect 1338 4655 1339 4659
rect 1344 4655 1345 4659
rect 1350 4655 1351 4659
rect 1356 4655 1357 4659
rect 1362 4655 1363 4659
rect 1744 4655 1745 4659
rect 1750 4655 1751 4659
rect 1756 4655 1757 4659
rect 1762 4655 1763 4659
rect 1768 4655 1769 4659
rect 1774 4655 1775 4659
rect 1019 4612 1020 4616
rect 1025 4612 1026 4616
rect 1031 4612 1032 4616
rect 1037 4612 1038 4616
rect 1043 4612 1044 4616
rect 1049 4612 1050 4616
rect 1109 4612 1110 4616
rect 1115 4612 1116 4616
rect 1121 4612 1122 4616
rect 1127 4612 1128 4616
rect 1133 4612 1134 4616
rect 1139 4612 1140 4616
rect 1493 4612 1494 4616
rect 1499 4612 1500 4616
rect 1505 4612 1506 4616
rect 1511 4612 1512 4616
rect 1517 4612 1518 4616
rect 1523 4612 1524 4616
rect 1583 4612 1584 4616
rect 1589 4612 1590 4616
rect 1595 4612 1596 4616
rect 1601 4612 1602 4616
rect 1607 4612 1608 4616
rect 1613 4612 1614 4616
rect 1967 4612 1968 4616
rect 1973 4612 1974 4616
rect 1979 4612 1980 4616
rect 1985 4612 1986 4616
rect 1991 4612 1992 4616
rect 1997 4612 1998 4616
rect 2057 4612 2058 4616
rect 2063 4612 2064 4616
rect 2069 4612 2070 4616
rect 2075 4612 2076 4616
rect 2081 4612 2082 4616
rect 2087 4612 2088 4616
rect 2915 4612 2916 4616
rect 2921 4612 2922 4616
rect 2927 4612 2928 4616
rect 2933 4612 2934 4616
rect 2939 4612 2940 4616
rect 2945 4612 2946 4616
rect 3005 4612 3006 4616
rect 3011 4612 3012 4616
rect 3017 4612 3018 4616
rect 3023 4612 3024 4616
rect 3029 4612 3030 4616
rect 3035 4612 3036 4616
rect 1019 4599 1020 4603
rect 1025 4599 1026 4603
rect 1031 4599 1032 4603
rect 1037 4599 1038 4603
rect 1043 4599 1044 4603
rect 1049 4599 1050 4603
rect 1109 4599 1110 4603
rect 1115 4599 1116 4603
rect 1121 4599 1122 4603
rect 1127 4599 1128 4603
rect 1133 4599 1134 4603
rect 1139 4599 1140 4603
rect 1493 4599 1494 4603
rect 1499 4599 1500 4603
rect 1505 4599 1506 4603
rect 1511 4599 1512 4603
rect 1517 4599 1518 4603
rect 1523 4599 1524 4603
rect 1583 4599 1584 4603
rect 1589 4599 1590 4603
rect 1595 4599 1596 4603
rect 1601 4599 1602 4603
rect 1607 4599 1608 4603
rect 1613 4599 1614 4603
rect 1967 4599 1968 4603
rect 1973 4599 1974 4603
rect 1979 4599 1980 4603
rect 1985 4599 1986 4603
rect 1991 4599 1992 4603
rect 1997 4599 1998 4603
rect 2057 4599 2058 4603
rect 2063 4599 2064 4603
rect 2069 4599 2070 4603
rect 2075 4599 2076 4603
rect 2081 4599 2082 4603
rect 2087 4599 2088 4603
rect 2915 4599 2916 4603
rect 2921 4599 2922 4603
rect 2927 4599 2928 4603
rect 2933 4599 2934 4603
rect 2939 4599 2940 4603
rect 2945 4599 2946 4603
rect 3005 4599 3006 4603
rect 3011 4599 3012 4603
rect 3017 4599 3018 4603
rect 3023 4599 3024 4603
rect 3029 4599 3030 4603
rect 3035 4599 3036 4603
rect 1020 4583 1021 4586
rect 1026 4583 1027 4586
rect 1032 4583 1033 4586
rect 1038 4583 1039 4586
rect 1120 4583 1121 4586
rect 1126 4583 1127 4586
rect 1132 4583 1133 4586
rect 1138 4583 1139 4586
rect 1494 4583 1495 4586
rect 1500 4583 1501 4586
rect 1506 4583 1507 4586
rect 1512 4583 1513 4586
rect 1594 4583 1595 4586
rect 1600 4583 1601 4586
rect 1606 4583 1607 4586
rect 1612 4583 1613 4586
rect 1968 4583 1969 4586
rect 1974 4583 1975 4586
rect 1980 4583 1981 4586
rect 1986 4583 1987 4586
rect 2068 4583 2069 4586
rect 2074 4583 2075 4586
rect 2080 4583 2081 4586
rect 2086 4583 2087 4586
rect 2916 4583 2917 4586
rect 2922 4583 2923 4586
rect 2928 4583 2929 4586
rect 2934 4583 2935 4586
rect 3016 4583 3017 4586
rect 3022 4583 3023 4586
rect 3028 4583 3029 4586
rect 3034 4583 3035 4586
rect 1014 4582 1018 4583
rect 1020 4582 1024 4583
rect 1026 4582 1030 4583
rect 1032 4582 1036 4583
rect 1038 4582 1042 4583
rect 1114 4582 1118 4583
rect 1120 4582 1124 4583
rect 1126 4582 1130 4583
rect 1132 4582 1136 4583
rect 1138 4582 1142 4583
rect 1488 4582 1492 4583
rect 1494 4582 1498 4583
rect 1500 4582 1504 4583
rect 1506 4582 1510 4583
rect 1512 4582 1516 4583
rect 1588 4582 1592 4583
rect 1594 4582 1598 4583
rect 1600 4582 1604 4583
rect 1606 4582 1610 4583
rect 1612 4582 1616 4583
rect 1962 4582 1966 4583
rect 1968 4582 1972 4583
rect 1974 4582 1978 4583
rect 1980 4582 1984 4583
rect 1986 4582 1990 4583
rect 2062 4582 2066 4583
rect 2068 4582 2072 4583
rect 2074 4582 2078 4583
rect 2080 4582 2084 4583
rect 2086 4582 2090 4583
rect 2910 4582 2914 4583
rect 2916 4582 2920 4583
rect 2922 4582 2926 4583
rect 2928 4582 2932 4583
rect 2934 4582 2938 4583
rect 3010 4582 3014 4583
rect 3016 4582 3020 4583
rect 3022 4582 3026 4583
rect 3028 4582 3032 4583
rect 3034 4582 3038 4583
rect 1020 4576 1021 4580
rect 1026 4576 1027 4580
rect 1032 4576 1033 4580
rect 1038 4576 1039 4580
rect 1120 4576 1121 4580
rect 1126 4576 1127 4580
rect 1132 4576 1133 4580
rect 1138 4576 1139 4580
rect 1494 4576 1495 4580
rect 1500 4576 1501 4580
rect 1506 4576 1507 4580
rect 1512 4576 1513 4580
rect 1594 4576 1595 4580
rect 1600 4576 1601 4580
rect 1606 4576 1607 4580
rect 1612 4576 1613 4580
rect 1968 4576 1969 4580
rect 1974 4576 1975 4580
rect 1980 4576 1981 4580
rect 1986 4576 1987 4580
rect 2068 4576 2069 4580
rect 2074 4576 2075 4580
rect 2080 4576 2081 4580
rect 2086 4576 2087 4580
rect 2916 4576 2917 4580
rect 2922 4576 2923 4580
rect 2928 4576 2929 4580
rect 2934 4576 2935 4580
rect 3016 4576 3017 4580
rect 3022 4576 3023 4580
rect 3028 4576 3029 4580
rect 3034 4576 3035 4580
rect 1020 4570 1021 4573
rect 1026 4570 1027 4573
rect 1032 4570 1033 4573
rect 1038 4570 1039 4573
rect 1120 4570 1121 4573
rect 1126 4570 1127 4573
rect 1132 4570 1133 4573
rect 1138 4570 1139 4573
rect 1494 4570 1495 4573
rect 1500 4570 1501 4573
rect 1506 4570 1507 4573
rect 1512 4570 1513 4573
rect 1594 4570 1595 4573
rect 1600 4570 1601 4573
rect 1606 4570 1607 4573
rect 1612 4570 1613 4573
rect 1968 4570 1969 4573
rect 1974 4570 1975 4573
rect 1980 4570 1981 4573
rect 1986 4570 1987 4573
rect 2068 4570 2069 4573
rect 2074 4570 2075 4573
rect 2080 4570 2081 4573
rect 2086 4570 2087 4573
rect 2916 4570 2917 4573
rect 2922 4570 2923 4573
rect 2928 4570 2929 4573
rect 2934 4570 2935 4573
rect 3016 4570 3017 4573
rect 3022 4570 3023 4573
rect 3028 4570 3029 4573
rect 3034 4570 3035 4573
rect 1014 4569 1018 4570
rect 1020 4569 1024 4570
rect 1026 4569 1030 4570
rect 1032 4569 1036 4570
rect 1038 4569 1042 4570
rect 1114 4569 1118 4570
rect 1120 4569 1124 4570
rect 1126 4569 1130 4570
rect 1132 4569 1136 4570
rect 1138 4569 1142 4570
rect 1488 4569 1492 4570
rect 1494 4569 1498 4570
rect 1500 4569 1504 4570
rect 1506 4569 1510 4570
rect 1512 4569 1516 4570
rect 1588 4569 1592 4570
rect 1594 4569 1598 4570
rect 1600 4569 1604 4570
rect 1606 4569 1610 4570
rect 1612 4569 1616 4570
rect 1962 4569 1966 4570
rect 1968 4569 1972 4570
rect 1974 4569 1978 4570
rect 1980 4569 1984 4570
rect 1986 4569 1990 4570
rect 2062 4569 2066 4570
rect 2068 4569 2072 4570
rect 2074 4569 2078 4570
rect 2080 4569 2084 4570
rect 2086 4569 2090 4570
rect 2910 4569 2914 4570
rect 2916 4569 2920 4570
rect 2922 4569 2926 4570
rect 2928 4569 2932 4570
rect 2934 4569 2938 4570
rect 3010 4569 3014 4570
rect 3016 4569 3020 4570
rect 3022 4569 3026 4570
rect 3028 4569 3032 4570
rect 3034 4569 3038 4570
rect 1020 4564 1021 4567
rect 1026 4564 1027 4567
rect 1032 4564 1033 4567
rect 1038 4564 1039 4567
rect 1120 4564 1121 4567
rect 1126 4564 1127 4567
rect 1132 4564 1133 4567
rect 1138 4564 1139 4567
rect 1494 4564 1495 4567
rect 1500 4564 1501 4567
rect 1506 4564 1507 4567
rect 1512 4564 1513 4567
rect 1594 4564 1595 4567
rect 1600 4564 1601 4567
rect 1606 4564 1607 4567
rect 1612 4564 1613 4567
rect 1968 4564 1969 4567
rect 1974 4564 1975 4567
rect 1980 4564 1981 4567
rect 1986 4564 1987 4567
rect 2068 4564 2069 4567
rect 2074 4564 2075 4567
rect 2080 4564 2081 4567
rect 2086 4564 2087 4567
rect 2916 4564 2917 4567
rect 2922 4564 2923 4567
rect 2928 4564 2929 4567
rect 2934 4564 2935 4567
rect 3016 4564 3017 4567
rect 3022 4564 3023 4567
rect 3028 4564 3029 4567
rect 3034 4564 3035 4567
rect 1014 4563 1018 4564
rect 1020 4563 1024 4564
rect 1026 4563 1030 4564
rect 1032 4563 1036 4564
rect 1038 4563 1042 4564
rect 1114 4563 1118 4564
rect 1120 4563 1124 4564
rect 1126 4563 1130 4564
rect 1132 4563 1136 4564
rect 1138 4563 1142 4564
rect 1488 4563 1492 4564
rect 1494 4563 1498 4564
rect 1500 4563 1504 4564
rect 1506 4563 1510 4564
rect 1512 4563 1516 4564
rect 1588 4563 1592 4564
rect 1594 4563 1598 4564
rect 1600 4563 1604 4564
rect 1606 4563 1610 4564
rect 1612 4563 1616 4564
rect 1962 4563 1966 4564
rect 1968 4563 1972 4564
rect 1974 4563 1978 4564
rect 1980 4563 1984 4564
rect 1986 4563 1990 4564
rect 2062 4563 2066 4564
rect 2068 4563 2072 4564
rect 2074 4563 2078 4564
rect 2080 4563 2084 4564
rect 2086 4563 2090 4564
rect 2910 4563 2914 4564
rect 2916 4563 2920 4564
rect 2922 4563 2926 4564
rect 2928 4563 2932 4564
rect 2934 4563 2938 4564
rect 3010 4563 3014 4564
rect 3016 4563 3020 4564
rect 3022 4563 3026 4564
rect 3028 4563 3032 4564
rect 3034 4563 3038 4564
rect 1020 4558 1021 4561
rect 1026 4558 1027 4561
rect 1032 4558 1033 4561
rect 1038 4558 1039 4561
rect 1120 4558 1121 4561
rect 1126 4558 1127 4561
rect 1132 4558 1133 4561
rect 1138 4558 1139 4561
rect 1494 4558 1495 4561
rect 1500 4558 1501 4561
rect 1506 4558 1507 4561
rect 1512 4558 1513 4561
rect 1594 4558 1595 4561
rect 1600 4558 1601 4561
rect 1606 4558 1607 4561
rect 1612 4558 1613 4561
rect 1968 4558 1969 4561
rect 1974 4558 1975 4561
rect 1980 4558 1981 4561
rect 1986 4558 1987 4561
rect 2068 4558 2069 4561
rect 2074 4558 2075 4561
rect 2080 4558 2081 4561
rect 2086 4558 2087 4561
rect 2916 4558 2917 4561
rect 2922 4558 2923 4561
rect 2928 4558 2929 4561
rect 2934 4558 2935 4561
rect 3016 4558 3017 4561
rect 3022 4558 3023 4561
rect 3028 4558 3029 4561
rect 3034 4558 3035 4561
rect 1014 4557 1018 4558
rect 1020 4557 1024 4558
rect 1026 4557 1030 4558
rect 1032 4557 1036 4558
rect 1038 4557 1042 4558
rect 1114 4557 1118 4558
rect 1120 4557 1124 4558
rect 1126 4557 1130 4558
rect 1132 4557 1136 4558
rect 1138 4557 1142 4558
rect 1488 4557 1492 4558
rect 1494 4557 1498 4558
rect 1500 4557 1504 4558
rect 1506 4557 1510 4558
rect 1512 4557 1516 4558
rect 1588 4557 1592 4558
rect 1594 4557 1598 4558
rect 1600 4557 1604 4558
rect 1606 4557 1610 4558
rect 1612 4557 1616 4558
rect 1962 4557 1966 4558
rect 1968 4557 1972 4558
rect 1974 4557 1978 4558
rect 1980 4557 1984 4558
rect 1986 4557 1990 4558
rect 2062 4557 2066 4558
rect 2068 4557 2072 4558
rect 2074 4557 2078 4558
rect 2080 4557 2084 4558
rect 2086 4557 2090 4558
rect 2910 4557 2914 4558
rect 2916 4557 2920 4558
rect 2922 4557 2926 4558
rect 2928 4557 2932 4558
rect 2934 4557 2938 4558
rect 3010 4557 3014 4558
rect 3016 4557 3020 4558
rect 3022 4557 3026 4558
rect 3028 4557 3032 4558
rect 3034 4557 3038 4558
rect 1020 4551 1021 4555
rect 1026 4551 1027 4555
rect 1032 4551 1033 4555
rect 1038 4551 1039 4555
rect 1120 4551 1121 4555
rect 1126 4551 1127 4555
rect 1132 4551 1133 4555
rect 1138 4551 1139 4555
rect 1494 4551 1495 4555
rect 1500 4551 1501 4555
rect 1506 4551 1507 4555
rect 1512 4551 1513 4555
rect 1594 4551 1595 4555
rect 1600 4551 1601 4555
rect 1606 4551 1607 4555
rect 1612 4551 1613 4555
rect 1968 4551 1969 4555
rect 1974 4551 1975 4555
rect 1980 4551 1981 4555
rect 1986 4551 1987 4555
rect 2068 4551 2069 4555
rect 2074 4551 2075 4555
rect 2080 4551 2081 4555
rect 2086 4551 2087 4555
rect 2916 4551 2917 4555
rect 2922 4551 2923 4555
rect 2928 4551 2929 4555
rect 2934 4551 2935 4555
rect 3016 4551 3017 4555
rect 3022 4551 3023 4555
rect 3028 4551 3029 4555
rect 3034 4551 3035 4555
rect 1019 4525 1020 4529
rect 1025 4525 1026 4529
rect 1031 4525 1032 4529
rect 1037 4525 1038 4529
rect 1043 4525 1044 4529
rect 1049 4525 1050 4529
rect 1109 4525 1110 4529
rect 1115 4525 1116 4529
rect 1121 4525 1122 4529
rect 1127 4525 1128 4529
rect 1133 4525 1134 4529
rect 1139 4525 1140 4529
rect 1493 4525 1494 4529
rect 1499 4525 1500 4529
rect 1505 4525 1506 4529
rect 1511 4525 1512 4529
rect 1517 4525 1518 4529
rect 1523 4525 1524 4529
rect 1583 4525 1584 4529
rect 1589 4525 1590 4529
rect 1595 4525 1596 4529
rect 1601 4525 1602 4529
rect 1607 4525 1608 4529
rect 1613 4525 1614 4529
rect 1967 4525 1968 4529
rect 1973 4525 1974 4529
rect 1979 4525 1980 4529
rect 1985 4525 1986 4529
rect 1991 4525 1992 4529
rect 1997 4525 1998 4529
rect 2057 4525 2058 4529
rect 2063 4525 2064 4529
rect 2069 4525 2070 4529
rect 2075 4525 2076 4529
rect 2081 4525 2082 4529
rect 2087 4525 2088 4529
rect 2915 4525 2916 4529
rect 2921 4525 2922 4529
rect 2927 4525 2928 4529
rect 2933 4525 2934 4529
rect 2939 4525 2940 4529
rect 2945 4525 2946 4529
rect 3005 4525 3006 4529
rect 3011 4525 3012 4529
rect 3017 4525 3018 4529
rect 3023 4525 3024 4529
rect 3029 4525 3030 4529
rect 3035 4525 3036 4529
rect 1019 4507 1020 4511
rect 1025 4507 1026 4511
rect 1031 4507 1032 4511
rect 1037 4507 1038 4511
rect 1043 4507 1044 4511
rect 1049 4507 1050 4511
rect 1109 4507 1110 4511
rect 1115 4507 1116 4511
rect 1121 4507 1122 4511
rect 1127 4507 1128 4511
rect 1133 4507 1134 4511
rect 1139 4507 1140 4511
rect 1493 4507 1494 4511
rect 1499 4507 1500 4511
rect 1505 4507 1506 4511
rect 1511 4507 1512 4511
rect 1517 4507 1518 4511
rect 1523 4507 1524 4511
rect 1583 4507 1584 4511
rect 1589 4507 1590 4511
rect 1595 4507 1596 4511
rect 1601 4507 1602 4511
rect 1607 4507 1608 4511
rect 1613 4507 1614 4511
rect 1967 4507 1968 4511
rect 1973 4507 1974 4511
rect 1979 4507 1980 4511
rect 1985 4507 1986 4511
rect 1991 4507 1992 4511
rect 1997 4507 1998 4511
rect 2057 4507 2058 4511
rect 2063 4507 2064 4511
rect 2069 4507 2070 4511
rect 2075 4507 2076 4511
rect 2081 4507 2082 4511
rect 2087 4507 2088 4511
rect 2915 4507 2916 4511
rect 2921 4507 2922 4511
rect 2927 4507 2928 4511
rect 2933 4507 2934 4511
rect 2939 4507 2940 4511
rect 2945 4507 2946 4511
rect 3005 4507 3006 4511
rect 3011 4507 3012 4511
rect 3017 4507 3018 4511
rect 3023 4507 3024 4511
rect 3029 4507 3030 4511
rect 3035 4507 3036 4511
rect 3665 4203 3671 4206
rect 3695 4196 3707 4197
rect 3699 4192 3703 4193
<< nwell >>
rect 3370 4228 3515 4378
<< ptransistor >>
rect 3398 4245 3404 4365
rect 3419 4245 3425 4365
rect 3440 4245 3446 4365
<< pdiffusion >>
rect 3392 4364 3398 4365
rect 3392 4290 3393 4364
rect 3397 4290 3398 4364
rect 3392 4268 3398 4290
rect 3392 4246 3393 4268
rect 3397 4246 3398 4268
rect 3392 4245 3398 4246
rect 3404 4364 3410 4365
rect 3404 4358 3405 4364
rect 3409 4358 3410 4364
rect 3404 4354 3410 4358
rect 3404 4350 3405 4354
rect 3409 4350 3410 4354
rect 3404 4346 3410 4350
rect 3404 4342 3405 4346
rect 3409 4342 3410 4346
rect 3404 4338 3410 4342
rect 3404 4334 3405 4338
rect 3409 4334 3410 4338
rect 3404 4330 3410 4334
rect 3404 4326 3405 4330
rect 3409 4326 3410 4330
rect 3404 4322 3410 4326
rect 3404 4318 3405 4322
rect 3409 4318 3410 4322
rect 3404 4314 3410 4318
rect 3404 4310 3405 4314
rect 3409 4310 3410 4314
rect 3404 4306 3410 4310
rect 3404 4302 3405 4306
rect 3409 4302 3410 4306
rect 3404 4298 3410 4302
rect 3404 4294 3405 4298
rect 3409 4294 3410 4298
rect 3404 4290 3410 4294
rect 3404 4286 3405 4290
rect 3409 4286 3410 4290
rect 3404 4282 3410 4286
rect 3404 4278 3405 4282
rect 3409 4278 3410 4282
rect 3404 4274 3410 4278
rect 3404 4270 3405 4274
rect 3409 4270 3410 4274
rect 3404 4266 3410 4270
rect 3404 4262 3405 4266
rect 3409 4262 3410 4266
rect 3404 4258 3410 4262
rect 3404 4254 3405 4258
rect 3409 4254 3410 4258
rect 3404 4250 3410 4254
rect 3404 4246 3405 4250
rect 3409 4246 3410 4250
rect 3404 4245 3410 4246
rect 3413 4364 3419 4365
rect 3413 4246 3414 4364
rect 3418 4246 3419 4364
rect 3413 4245 3419 4246
rect 3425 4364 3431 4365
rect 3425 4358 3426 4364
rect 3430 4358 3431 4364
rect 3425 4354 3431 4358
rect 3425 4350 3426 4354
rect 3430 4350 3431 4354
rect 3425 4346 3431 4350
rect 3425 4342 3426 4346
rect 3430 4342 3431 4346
rect 3425 4338 3431 4342
rect 3425 4334 3426 4338
rect 3430 4334 3431 4338
rect 3425 4330 3431 4334
rect 3425 4326 3426 4330
rect 3430 4326 3431 4330
rect 3425 4322 3431 4326
rect 3425 4318 3426 4322
rect 3430 4318 3431 4322
rect 3425 4314 3431 4318
rect 3425 4310 3426 4314
rect 3430 4310 3431 4314
rect 3425 4306 3431 4310
rect 3425 4302 3426 4306
rect 3430 4302 3431 4306
rect 3425 4298 3431 4302
rect 3425 4294 3426 4298
rect 3430 4294 3431 4298
rect 3425 4290 3431 4294
rect 3425 4286 3426 4290
rect 3430 4286 3431 4290
rect 3425 4282 3431 4286
rect 3425 4278 3426 4282
rect 3430 4278 3431 4282
rect 3425 4274 3431 4278
rect 3425 4270 3426 4274
rect 3430 4270 3431 4274
rect 3425 4266 3431 4270
rect 3425 4262 3426 4266
rect 3430 4262 3431 4266
rect 3425 4258 3431 4262
rect 3425 4254 3426 4258
rect 3430 4254 3431 4258
rect 3425 4250 3431 4254
rect 3425 4246 3426 4250
rect 3430 4246 3431 4250
rect 3425 4245 3431 4246
rect 3434 4364 3440 4365
rect 3434 4246 3435 4364
rect 3439 4246 3440 4364
rect 3434 4245 3440 4246
rect 3446 4364 3452 4365
rect 3446 4358 3447 4364
rect 3451 4358 3452 4364
rect 3446 4354 3452 4358
rect 3446 4350 3447 4354
rect 3451 4350 3452 4354
rect 3446 4346 3452 4350
rect 3446 4342 3447 4346
rect 3451 4342 3452 4346
rect 3446 4338 3452 4342
rect 3446 4334 3447 4338
rect 3451 4334 3452 4338
rect 3446 4330 3452 4334
rect 3446 4326 3447 4330
rect 3451 4326 3452 4330
rect 3446 4322 3452 4326
rect 3446 4318 3447 4322
rect 3451 4318 3452 4322
rect 3446 4314 3452 4318
rect 3446 4310 3447 4314
rect 3451 4310 3452 4314
rect 3446 4306 3452 4310
rect 3446 4302 3447 4306
rect 3451 4302 3452 4306
rect 3446 4298 3452 4302
rect 3446 4294 3447 4298
rect 3451 4294 3452 4298
rect 3446 4290 3452 4294
rect 3446 4286 3447 4290
rect 3451 4286 3452 4290
rect 3446 4282 3452 4286
rect 3446 4278 3447 4282
rect 3451 4278 3452 4282
rect 3446 4274 3452 4278
rect 3446 4270 3447 4274
rect 3451 4270 3452 4274
rect 3446 4266 3452 4270
rect 3446 4262 3447 4266
rect 3451 4262 3452 4266
rect 3446 4258 3452 4262
rect 3446 4254 3447 4258
rect 3451 4254 3452 4258
rect 3446 4250 3452 4254
rect 3446 4246 3447 4250
rect 3451 4246 3452 4250
rect 3446 4245 3452 4246
<< pdcontact >>
rect 3393 4290 3397 4364
rect 3393 4246 3397 4268
rect 3405 4358 3409 4364
rect 3405 4350 3409 4354
rect 3405 4342 3409 4346
rect 3405 4334 3409 4338
rect 3405 4326 3409 4330
rect 3405 4318 3409 4322
rect 3405 4310 3409 4314
rect 3405 4302 3409 4306
rect 3405 4294 3409 4298
rect 3405 4286 3409 4290
rect 3405 4278 3409 4282
rect 3405 4270 3409 4274
rect 3405 4262 3409 4266
rect 3405 4254 3409 4258
rect 3405 4246 3409 4250
rect 3414 4246 3418 4364
rect 3426 4358 3430 4364
rect 3426 4350 3430 4354
rect 3426 4342 3430 4346
rect 3426 4334 3430 4338
rect 3426 4326 3430 4330
rect 3426 4318 3430 4322
rect 3426 4310 3430 4314
rect 3426 4302 3430 4306
rect 3426 4294 3430 4298
rect 3426 4286 3430 4290
rect 3426 4278 3430 4282
rect 3426 4270 3430 4274
rect 3426 4262 3430 4266
rect 3426 4254 3430 4258
rect 3426 4246 3430 4250
rect 3435 4246 3439 4364
rect 3447 4358 3451 4364
rect 3447 4350 3451 4354
rect 3447 4342 3451 4346
rect 3447 4334 3451 4338
rect 3447 4326 3451 4330
rect 3447 4318 3451 4322
rect 3447 4310 3451 4314
rect 3447 4302 3451 4306
rect 3447 4294 3451 4298
rect 3447 4286 3451 4290
rect 3447 4278 3451 4282
rect 3447 4270 3451 4274
rect 3447 4262 3451 4266
rect 3447 4254 3451 4258
rect 3447 4246 3451 4250
<< nsubstratencontact >>
rect 3463 4250 3508 4358
<< polysilicon >>
rect 3215 4369 3221 4374
rect 3398 4372 3446 4373
rect 3398 4367 3399 4372
rect 3445 4367 3446 4372
rect 3398 4366 3446 4367
rect 3398 4365 3404 4366
rect 3419 4365 3425 4366
rect 3440 4365 3446 4366
rect 3808 4358 3814 4363
rect 3398 4244 3404 4245
rect 3419 4244 3425 4245
rect 3440 4244 3446 4245
rect 3398 4243 3446 4244
rect 3398 4238 3399 4243
rect 3430 4238 3446 4243
rect 3398 4237 3446 4238
<< polycontact >>
rect 3399 4367 3445 4372
rect 3399 4238 3430 4243
<< metal1 >>
rect 1182 4528 1244 4529
rect 1013 4390 1053 4496
rect 1070 4404 1086 4496
rect 1159 4487 1244 4528
rect 1175 4486 1244 4487
rect 1198 4452 1244 4486
rect 1544 4474 1560 4507
rect 2018 4482 2034 4504
rect 1250 4404 1560 4474
rect 2006 4473 2047 4482
rect 1070 4393 1096 4404
rect 1244 4400 1560 4404
rect 1244 4393 1731 4397
rect 1013 4272 1101 4390
rect 1252 4381 1731 4393
rect 1289 4375 1731 4381
rect 1289 4316 1737 4375
rect 1576 3948 1737 4316
rect 1981 4056 2072 4473
rect 2865 4067 2904 4500
rect 2910 4383 2948 4502
rect 3182 4463 3200 4464
rect 3182 4462 3346 4463
rect 3440 4462 3456 4511
rect 3182 4447 3456 4462
rect 3857 4460 3897 4489
rect 2910 4357 3176 4383
rect 3182 4364 3200 4447
rect 3344 4446 3456 4447
rect 3782 4418 3793 4419
rect 3782 4388 3784 4418
rect 3791 4388 3793 4418
rect 3414 4364 3418 4367
rect 2910 4343 3121 4357
rect 2910 4330 3058 4343
rect 3451 4358 3507 4359
rect 3451 4250 3463 4358
rect 3782 4354 3793 4388
rect 3817 4382 3897 4460
rect 3817 4346 3853 4382
rect 2865 4064 3051 4067
rect 1979 4007 2838 4056
rect 2865 4034 3214 4064
rect 3236 4007 3289 4246
rect 3414 4243 3418 4246
rect 3435 4242 3439 4246
rect 3435 4234 3458 4242
rect 3914 4238 3930 4505
rect 3431 4097 3458 4234
rect 3826 4236 3930 4238
rect 3826 4206 3897 4236
rect 3927 4206 3930 4236
rect 3826 4202 3930 4206
rect 3431 4095 3635 4097
rect 3431 4061 3638 4095
rect 3991 4090 4031 4494
rect 4049 4404 4135 4405
rect 4045 4388 4492 4404
rect 4045 4366 4467 4388
rect 3431 4060 3635 4061
rect 3771 4051 4031 4090
rect 1979 3962 3289 4007
rect 2769 3961 3289 3962
rect 1576 3947 3599 3948
rect 4049 3947 4134 4366
rect 1576 3847 4134 3947
rect 4209 3991 4491 4031
rect 4209 3830 4265 3991
rect 1437 3794 1515 3809
rect 1437 3788 3587 3794
rect 1437 3721 3546 3788
rect 3578 3721 3587 3788
rect 3973 3780 4265 3830
rect 4374 3914 4491 3930
rect 1437 3716 3587 3721
rect 1437 606 1515 3716
rect 3889 3682 3925 3684
rect 1561 3681 1562 3682
rect 3889 3681 3930 3682
rect 1556 3679 3930 3681
rect 1556 3585 3898 3679
rect 1556 3584 3925 3585
rect 1561 1075 1658 3584
rect 3889 3583 3925 3584
rect 3974 3527 4024 3780
rect 4374 3756 4452 3914
rect 4086 3663 4452 3756
rect 4089 3335 4158 3663
rect 4309 3440 4491 3456
rect 4013 3293 4158 3335
rect 4310 3212 4349 3440
rect 4014 3176 4349 3212
rect 4013 3054 4279 3089
rect 3699 3031 3770 3043
rect 3699 2871 3743 3031
rect 3752 2960 4215 3027
rect 4249 2982 4279 3054
rect 4249 2966 4491 2982
rect 3983 2959 4215 2960
rect 4158 2949 4215 2959
rect 4158 2909 4491 2949
rect 3699 2869 4311 2871
rect 3699 2864 4312 2869
rect 3700 2808 4312 2864
rect 4229 2526 4312 2808
rect 4229 2508 4483 2526
rect 4229 2492 4491 2508
rect 4229 2471 4483 2492
rect 4457 2034 4484 2037
rect 4457 2018 4490 2034
rect 4457 2017 4484 2018
rect 4447 1961 4490 2001
rect 1561 1064 1564 1075
rect 1655 1064 1658 1075
rect 1561 1061 1658 1064
rect 1070 547 1521 606
rect 1070 508 1086 547
rect 1544 531 1554 1056
rect 4388 596 4490 612
rect 1544 512 1557 531
rect 1574 524 1661 535
rect 1621 510 1661 524
rect 4388 510 4404 596
<< m2contact >>
rect 3784 4388 3791 4418
rect 3216 4368 3220 4372
rect 3393 4268 3397 4290
rect 3405 4354 3409 4358
rect 3405 4346 3409 4350
rect 3405 4338 3409 4342
rect 3405 4330 3409 4334
rect 3405 4322 3409 4326
rect 3405 4314 3409 4318
rect 3405 4306 3409 4310
rect 3405 4298 3409 4302
rect 3405 4290 3409 4294
rect 3405 4282 3409 4286
rect 3405 4274 3409 4278
rect 3405 4266 3409 4270
rect 3405 4258 3409 4262
rect 3405 4250 3409 4254
rect 3426 4354 3430 4358
rect 3426 4346 3430 4350
rect 3426 4338 3430 4342
rect 3426 4330 3430 4334
rect 3426 4322 3430 4326
rect 3426 4314 3430 4318
rect 3426 4306 3430 4310
rect 3426 4298 3430 4302
rect 3426 4290 3430 4294
rect 3426 4282 3430 4286
rect 3426 4274 3430 4278
rect 3426 4266 3430 4270
rect 3426 4258 3430 4262
rect 3426 4250 3430 4254
rect 3447 4354 3451 4358
rect 3447 4346 3451 4350
rect 3447 4338 3451 4342
rect 3447 4330 3451 4334
rect 3447 4322 3451 4326
rect 3447 4314 3451 4318
rect 3447 4306 3451 4310
rect 3447 4298 3451 4302
rect 3447 4290 3451 4294
rect 3447 4282 3451 4286
rect 3447 4274 3451 4278
rect 3447 4266 3451 4270
rect 3447 4258 3451 4262
rect 3447 4250 3451 4254
rect 3809 4358 3813 4362
rect 3040 4095 3044 4099
rect 3897 4206 3927 4236
rect 3546 3721 3578 3788
rect 3898 3585 3926 3679
rect 1564 1064 1655 1075
rect 1562 525 1569 561
<< metal2 >>
rect 3485 4491 3513 4492
rect 2492 4476 2508 4491
rect 2452 3560 2543 4476
rect 2966 4417 2982 4491
rect 2966 4400 3228 4417
rect 2966 4399 3037 4400
rect 3212 4372 3227 4400
rect 3212 4368 3216 4372
rect 3220 4368 3227 4372
rect 3212 4364 3227 4368
rect 3473 4364 3513 4491
rect 4388 4477 4404 4487
rect 3405 4358 3513 4364
rect 3409 4354 3426 4358
rect 3430 4354 3447 4358
rect 3451 4354 3513 4358
rect 3405 4350 3513 4354
rect 3409 4346 3426 4350
rect 3430 4346 3447 4350
rect 3451 4346 3513 4350
rect 3405 4342 3513 4346
rect 3409 4338 3426 4342
rect 3430 4338 3447 4342
rect 3451 4338 3513 4342
rect 3405 4334 3513 4338
rect 3409 4330 3426 4334
rect 3430 4330 3447 4334
rect 3451 4330 3513 4334
rect 3405 4326 3513 4330
rect 3409 4322 3426 4326
rect 3430 4322 3447 4326
rect 3451 4322 3513 4326
rect 3405 4318 3513 4322
rect 3409 4314 3426 4318
rect 3430 4314 3447 4318
rect 3451 4314 3513 4318
rect 3405 4310 3513 4314
rect 3409 4306 3426 4310
rect 3430 4306 3447 4310
rect 3451 4306 3513 4310
rect 3405 4302 3513 4306
rect 3409 4298 3426 4302
rect 3430 4298 3447 4302
rect 3451 4298 3513 4302
rect 3405 4294 3513 4298
rect 3106 4290 3395 4291
rect 3409 4290 3426 4294
rect 3430 4290 3447 4294
rect 3451 4290 3513 4294
rect 3106 4268 3393 4290
rect 3405 4286 3513 4290
rect 3409 4282 3426 4286
rect 3430 4282 3447 4286
rect 3451 4282 3513 4286
rect 3405 4278 3513 4282
rect 3409 4274 3426 4278
rect 3430 4274 3447 4278
rect 3451 4274 3513 4278
rect 3405 4270 3513 4274
rect 3106 4267 3395 4268
rect 3106 4266 3149 4267
rect 3409 4266 3426 4270
rect 3430 4266 3447 4270
rect 3451 4266 3513 4270
rect 3106 4172 3126 4266
rect 3405 4262 3513 4266
rect 3409 4258 3426 4262
rect 3430 4258 3447 4262
rect 3451 4258 3513 4262
rect 3405 4254 3513 4258
rect 3409 4250 3426 4254
rect 3430 4250 3447 4254
rect 3451 4250 3513 4254
rect 3405 4246 3513 4250
rect 3534 4419 3599 4420
rect 3534 4418 3793 4419
rect 3534 4388 3784 4418
rect 3791 4388 3793 4418
rect 3534 4387 3793 4388
rect 3039 4159 3126 4172
rect 3039 4099 3056 4159
rect 3039 4095 3040 4099
rect 3044 4095 3056 4099
rect 3039 4092 3056 4095
rect 3534 3788 3599 4387
rect 3805 4366 4404 4477
rect 3805 4362 3816 4366
rect 3805 4358 3809 4362
rect 3813 4358 3816 4362
rect 3805 4354 3816 4358
rect 3898 4236 3930 4246
rect 3927 4206 3930 4236
rect 3534 3721 3546 3788
rect 3578 3721 3599 3788
rect 3534 3714 3599 3721
rect 3898 3876 3930 4206
rect 3898 3679 3931 3876
rect 3926 3586 3931 3679
rect 2452 3513 3738 3560
rect 2452 3478 3782 3513
rect 2452 3477 3738 3478
rect 2452 3476 2543 3477
rect 1561 1075 1658 1080
rect 1561 1064 1564 1075
rect 1655 1064 1658 1075
rect 1561 561 1658 1064
rect 1561 525 1562 561
rect 1569 525 1658 561
rect 1561 524 1658 525
use blankpad  blankpad_11
timestamp 1259953556
transform -1 0 841 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_0
timestamp 1259953556
transform -1 0 1315 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_1
timestamp 1259953556
transform -1 0 1789 0 -1 5000
box -2 0 476 513
use inpad  inpad_9
timestamp 1259953556
transform -1 0 2263 0 -1 5000
box -2 0 476 513
use inpad  inpad_8
timestamp 1259953556
transform -1 0 2737 0 -1 5000
box -2 0 476 513
use inpad  inpad_7
timestamp 1259953556
transform -1 0 3211 0 -1 5000
box -2 0 476 513
use inpad  inpad_6
timestamp 1259953556
transform -1 0 3685 0 -1 5000
box -2 0 476 513
use inpad  inpad_5
timestamp 1259953556
transform -1 0 4159 0 -1 5000
box -2 0 476 513
use inpadp2  inpadp2_0
timestamp 1418813110
transform -1 0 4633 0 -1 5000
box -2 0 476 513
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 4487
box 0 0 5000 513
use 2-OR  2-OR_0
timestamp 1418434502
transform -1 0 1392 0 -1 4250
box 147 -223 302 -14
use blankpad  blankpad_27
timestamp 1259953556
transform 0 1 0 -1 0 4633
box -2 0 476 513
use Opamp  Opamp_0
timestamp 1418333453
transform 1 0 3221 0 1 4072
box -193 -11 77 303
use Opamp  Opamp_1
timestamp 1418333453
transform 1 0 3814 0 1 4062
box -193 -11 77 303
use inpad  inpad_3
timestamp 1259953556
transform 0 -1 5000 1 0 4159
box -2 0 476 513
use inpad  inpad_12
timestamp 1259953556
transform 0 1 0 -1 0 4159
box -2 0 476 513
use inpad  inpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 3685
box -2 0 476 513
use inpad  inpad_13
timestamp 1259953556
transform 0 1 0 -1 0 3685
box -2 0 476 513
use DAC  DAC_0
timestamp 1418788810
transform -1 0 4009 0 -1 3535
box -14 4 257 511
use inpad  inpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 3211
box -2 0 476 513
use inpad  inpad_14
timestamp 1259953556
transform 0 1 0 -1 0 3211
box -2 0 476 513
use inpad  inpad_15
timestamp 1259953556
transform 0 1 0 -1 0 2737
box -2 0 476 513
use inpad  inpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 2737
box -2 0 476 513
use inpad  inpad_11
timestamp 1259953556
transform 0 -1 5000 1 0 2263
box -2 0 476 513
use 50K_resistor  50K_resistor_0
timestamp 1418811347
transform -1 0 4601 0 -1 2225
box 143 188 207 270
use inpad  inpad_16
timestamp 1259953556
transform 0 1 0 -1 0 2263
box -2 0 476 513
use inpad  inpad_17
timestamp 1259953556
transform 0 1 0 -1 0 1789
box -2 0 476 513
use inpad  inpad_19
timestamp 1259953556
transform 0 -1 5000 1 0 1789
box -2 0 476 513
use blankpad  blankpad_8
timestamp 1259953556
transform 0 -1 5000 1 0 1315
box -2 0 476 513
use inpad  inpad_18
timestamp 1259953556
transform 0 1 0 -1 0 1315
box -2 0 476 513
use 2_200K_resistors  2_200K_resistors_0
timestamp 1418810336
transform 0 -1 1838 1 0 354
box 170 181 703 290
use blankpad  blankpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 841
box -2 0 476 513
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 367
box 2 2 513 4264
use blankpad  blankpad_29
timestamp 1259953556
transform 0 1 0 -1 0 841
box -2 0 476 513
use blankpad  blankpad_18
timestamp 1259953556
transform 1 0 367 0 1 0
box -2 0 476 513
use inpad  inpad_10
timestamp 1259953556
transform 1 0 841 0 1 0
box -2 0 476 513
use inpad  inpad_4
timestamp 1259953556
transform 1 0 1315 0 1 0
box -2 0 476 513
use blankpad  blankpad_25
timestamp 1259953556
transform 1 0 1789 0 1 0
box -2 0 476 513
use blankpad  blankpad_24
timestamp 1259953556
transform 1 0 2263 0 1 0
box -2 0 476 513
use blankpad  blankpad_23
timestamp 1259953556
transform 1 0 2737 0 1 0
box -2 0 476 513
use blankpad  blankpad_22
timestamp 1259953556
transform 1 0 3211 0 1 0
box -2 0 476 513
use blankpad  blankpad_21
timestamp 1259953556
transform 1 0 3685 0 1 0
box -2 0 476 513
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 4487 0 1 367
box 0 2 511 4264
use barepad  barepad_0
timestamp 1259953556
transform 0 -1 5000 1 0 367
box -2 0 476 513
use barepad  barepad_1
timestamp 1259953556
transform 1 0 4159 0 1 0
box -2 0 476 513
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 5000 513
<< end >>
