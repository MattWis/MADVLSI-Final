magic
tech scmos
timestamp 1418810336
<< electrode >>
rect 189 254 194 256
rect 202 254 207 256
rect 215 254 220 256
rect 228 254 233 256
rect 241 254 246 256
rect 254 254 259 256
rect 267 254 272 256
rect 280 254 285 256
rect 293 254 298 256
rect 306 254 311 256
rect 319 254 324 256
rect 332 254 337 256
rect 345 254 350 256
rect 358 254 363 256
rect 371 254 376 256
rect 384 254 389 256
rect 397 254 402 256
rect 410 254 415 256
rect 423 254 428 256
rect 436 254 441 256
rect 449 254 454 256
rect 462 254 467 256
rect 475 254 480 256
rect 488 254 493 256
rect 501 254 506 256
rect 514 254 519 256
rect 527 254 532 256
rect 540 254 545 256
rect 553 254 558 256
rect 566 254 571 256
rect 579 254 584 256
rect 592 254 597 256
rect 605 254 610 256
rect 618 254 623 256
rect 631 254 636 256
rect 644 254 649 256
rect 657 254 662 256
rect 670 254 675 256
rect 683 254 688 256
rect 696 254 701 256
rect 189 202 194 204
rect 202 202 207 204
rect 215 202 220 204
rect 228 202 233 204
rect 241 202 246 204
rect 254 202 259 204
rect 267 202 272 204
rect 280 202 285 204
rect 293 202 298 204
rect 306 202 311 204
rect 319 202 324 204
rect 332 202 337 204
rect 345 202 350 204
rect 358 202 363 204
rect 371 202 376 204
rect 384 202 389 204
rect 397 202 402 204
rect 410 202 415 204
rect 423 202 428 204
rect 436 202 441 204
rect 449 202 454 204
rect 462 202 467 204
rect 475 202 480 204
rect 488 202 493 204
rect 501 202 506 204
rect 514 202 519 204
rect 527 202 532 204
rect 540 202 545 204
rect 553 202 558 204
rect 566 202 571 204
rect 579 202 584 204
rect 592 202 597 204
rect 605 202 610 204
rect 618 202 623 204
rect 631 202 636 204
rect 644 202 649 204
rect 657 202 662 204
rect 670 202 675 204
rect 683 202 688 204
rect 696 202 701 204
<< genericpoly2contact >>
rect 189 256 194 263
rect 202 256 207 263
rect 215 256 220 263
rect 228 256 233 263
rect 241 256 246 263
rect 254 256 259 263
rect 267 256 272 263
rect 280 256 285 263
rect 293 256 298 263
rect 306 256 311 263
rect 319 256 324 263
rect 332 256 337 263
rect 345 256 350 263
rect 358 256 363 263
rect 371 256 376 263
rect 384 256 389 263
rect 397 256 402 263
rect 410 256 415 263
rect 423 256 428 263
rect 436 256 441 263
rect 449 256 454 263
rect 462 256 467 263
rect 475 256 480 263
rect 488 256 493 263
rect 501 256 506 263
rect 514 256 519 263
rect 527 256 532 263
rect 540 256 545 263
rect 553 256 558 263
rect 566 256 571 263
rect 579 256 584 263
rect 592 256 597 263
rect 605 256 610 263
rect 618 256 623 263
rect 631 256 636 263
rect 644 256 649 263
rect 657 256 662 263
rect 670 256 675 263
rect 683 256 688 263
rect 696 256 701 263
rect 189 195 194 202
rect 202 195 207 202
rect 215 195 220 202
rect 228 195 233 202
rect 241 195 246 202
rect 254 195 259 202
rect 267 195 272 202
rect 280 195 285 202
rect 293 195 298 202
rect 306 195 311 202
rect 319 195 324 202
rect 332 195 337 202
rect 345 195 350 202
rect 358 195 363 202
rect 371 195 376 202
rect 384 195 389 202
rect 397 195 402 202
rect 410 195 415 202
rect 423 195 428 202
rect 436 195 441 202
rect 449 195 454 202
rect 462 195 467 202
rect 475 195 480 202
rect 488 195 493 202
rect 501 195 506 202
rect 514 195 519 202
rect 527 195 532 202
rect 540 195 545 202
rect 553 195 558 202
rect 566 195 571 202
rect 579 195 584 202
rect 592 195 597 202
rect 605 195 610 202
rect 618 195 623 202
rect 631 195 636 202
rect 644 195 649 202
rect 657 195 662 202
rect 670 195 675 202
rect 683 195 688 202
rect 696 195 701 202
<< metal1 >>
rect 170 281 702 290
rect 170 268 208 277
rect 170 255 195 264
rect 201 255 208 268
rect 214 270 247 277
rect 214 255 221 270
rect 227 249 234 264
rect 240 255 247 270
rect 266 270 299 277
rect 253 249 260 264
rect 266 255 273 270
rect 227 242 260 249
rect 279 249 286 264
rect 292 255 299 270
rect 318 270 351 277
rect 305 249 312 264
rect 318 255 325 270
rect 279 242 312 249
rect 331 249 338 264
rect 344 255 351 270
rect 370 270 403 277
rect 357 249 364 264
rect 370 255 377 270
rect 331 242 364 249
rect 383 249 390 264
rect 396 255 403 270
rect 422 270 455 277
rect 409 249 416 264
rect 422 255 429 270
rect 383 242 416 249
rect 435 249 442 264
rect 448 255 455 270
rect 474 270 507 277
rect 461 249 468 264
rect 474 255 481 270
rect 435 242 468 249
rect 487 249 494 264
rect 500 255 507 270
rect 526 270 559 277
rect 513 249 520 264
rect 526 255 533 270
rect 487 242 520 249
rect 539 249 546 264
rect 552 255 559 270
rect 578 270 611 277
rect 565 249 572 264
rect 578 255 585 270
rect 539 242 572 249
rect 591 249 598 264
rect 604 255 611 270
rect 630 270 663 277
rect 617 249 624 264
rect 630 255 637 270
rect 591 242 624 249
rect 643 249 650 264
rect 656 255 663 270
rect 669 249 676 264
rect 682 255 702 281
rect 643 242 676 249
rect 188 209 221 216
rect 188 194 195 209
rect 201 188 208 203
rect 214 194 221 209
rect 240 209 273 216
rect 227 188 234 203
rect 240 194 247 209
rect 201 181 234 188
rect 253 188 260 203
rect 266 194 273 209
rect 292 209 325 216
rect 279 188 286 203
rect 292 194 299 209
rect 253 181 286 188
rect 305 188 312 203
rect 318 194 325 209
rect 344 209 377 216
rect 331 188 338 203
rect 344 194 351 209
rect 305 181 338 188
rect 357 188 364 203
rect 370 194 377 209
rect 396 209 429 216
rect 383 188 390 203
rect 396 194 403 209
rect 357 181 390 188
rect 409 188 416 203
rect 422 194 429 209
rect 448 209 481 216
rect 435 188 442 203
rect 448 194 455 209
rect 409 181 442 188
rect 461 188 468 203
rect 474 194 481 209
rect 500 209 533 216
rect 487 188 494 203
rect 500 194 507 209
rect 461 181 494 188
rect 513 188 520 203
rect 526 194 533 209
rect 552 209 585 216
rect 539 188 546 203
rect 552 194 559 209
rect 513 181 546 188
rect 565 188 572 203
rect 578 194 585 209
rect 604 209 637 216
rect 591 188 598 203
rect 604 194 611 209
rect 565 181 598 188
rect 617 188 624 203
rect 630 194 637 209
rect 656 209 689 216
rect 643 188 650 203
rect 656 194 663 209
rect 617 181 650 188
rect 669 188 676 203
rect 682 194 689 209
rect 695 188 702 203
rect 669 181 702 188
<< high_resist >>
rect 187 204 189 254
rect 194 204 196 254
rect 200 204 202 254
rect 207 204 209 254
rect 213 204 215 254
rect 220 204 222 254
rect 226 204 228 254
rect 233 204 235 254
rect 239 204 241 254
rect 246 204 248 254
rect 252 204 254 254
rect 259 204 261 254
rect 265 204 267 254
rect 272 204 274 254
rect 278 204 280 254
rect 285 204 287 254
rect 291 204 293 254
rect 298 204 300 254
rect 304 204 306 254
rect 311 204 313 254
rect 317 204 319 254
rect 324 204 326 254
rect 330 204 332 254
rect 337 204 339 254
rect 343 204 345 254
rect 350 204 352 254
rect 356 204 358 254
rect 363 204 365 254
rect 369 204 371 254
rect 376 204 378 254
rect 382 204 384 254
rect 389 204 391 254
rect 395 204 397 254
rect 402 204 404 254
rect 408 204 410 254
rect 415 204 417 254
rect 421 204 423 254
rect 428 204 430 254
rect 434 204 436 254
rect 441 204 443 254
rect 447 204 449 254
rect 454 204 456 254
rect 460 204 462 254
rect 467 204 469 254
rect 473 204 475 254
rect 480 204 482 254
rect 486 204 488 254
rect 493 204 495 254
rect 499 204 501 254
rect 506 204 508 254
rect 512 204 514 254
rect 519 204 521 254
rect 525 204 527 254
rect 532 204 534 254
rect 538 204 540 254
rect 545 204 547 254
rect 551 204 553 254
rect 558 204 560 254
rect 564 204 566 254
rect 571 204 573 254
rect 577 204 579 254
rect 584 204 586 254
rect 590 204 592 254
rect 597 204 599 254
rect 603 204 605 254
rect 610 204 612 254
rect 616 204 618 254
rect 623 204 625 254
rect 629 204 631 254
rect 636 204 638 254
rect 642 204 644 254
rect 649 204 651 254
rect 655 204 657 254
rect 662 204 664 254
rect 668 204 670 254
rect 675 204 677 254
rect 681 204 683 254
rect 688 204 690 254
rect 694 204 696 254
rect 701 204 703 254
<< poly2_high_resist >>
rect 189 204 194 254
rect 202 204 207 254
rect 215 204 220 254
rect 228 204 233 254
rect 241 204 246 254
rect 254 204 259 254
rect 267 204 272 254
rect 280 204 285 254
rect 293 204 298 254
rect 306 204 311 254
rect 319 204 324 254
rect 332 204 337 254
rect 345 204 350 254
rect 358 204 363 254
rect 371 204 376 254
rect 384 204 389 254
rect 397 204 402 254
rect 410 204 415 254
rect 423 204 428 254
rect 436 204 441 254
rect 449 204 454 254
rect 462 204 467 254
rect 475 204 480 254
rect 488 204 493 254
rect 501 204 506 254
rect 514 204 519 254
rect 527 204 532 254
rect 540 204 545 254
rect 553 204 558 254
rect 566 204 571 254
rect 579 204 584 254
rect 592 204 597 254
rect 605 204 610 254
rect 618 204 623 254
rect 631 204 636 254
rect 644 204 649 254
rect 657 204 662 254
rect 670 204 675 254
rect 683 204 688 254
rect 696 204 701 254
<< end >>
