* SPICE3 file created from 2-OR.ext - technology: scmos

M1000 a_165_n141# B a_153_n141# w_147_n150# pfet w=1.8u l=0.6u
+  ad=1.62p pd=5.4u as=5.4p ps=9.6u
M1001 w_147_n150# A a_165_n141# w_147_n150# pfet w=1.8u l=0.6u
+  ad=459.54p pd=541.2u as=0p ps=0u
M1002 a_180_n144# a_153_n141# w_147_n150# w_147_n150# pfet w=3.6u l=0.6u
+  ad=6.48p pd=10.8u as=0p ps=0u
M1003 a_199_n216# a_180_n144# w_147_n150# w_147_n150# pfet w=36u l=0.6u
+  ad=64.8p pd=75.6u as=0p ps=0u
M1004 Z a_199_n216# w_147_n150# w_147_n150# pfet w=36u l=0.6u M=10
+  ad=324p pd=378u as=0p ps=0u
M1005 a_153_n141# B Gnd Gnd nfet w=1.8u l=0.6u
+  ad=6.48p pd=10.8u as=233.28p ps=291.6u
M1006 Gnd A a_153_n141# Gnd nfet w=1.8u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_180_n144# a_153_n141# Gnd Gnd nfet w=1.8u l=0.6u
+  ad=3.24p pd=7.2u as=0p ps=0u
M1008 a_199_n216# a_180_n144# Gnd Gnd nfet w=18u l=0.6u
+  ad=32.4p pd=39.6u as=0p ps=0u
M1009 Z a_199_n216# Gnd Gnd nfet w=18u l=0.6u M=10
+  ad=162p pd=198u as=0p ps=0u
