magic
tech scmos
timestamp 1418825699
<< m3contact >>
rect 1897 1889 1902 1894
rect 0 0 4 4
<< metal3 >>
rect 0 3795 3800 3800
rect 0 5 5 3795
rect -1 4 5 5
rect -1 0 0 4
rect 4 0 5 4
rect 8 3787 3792 3792
rect 8 5 13 3787
rect 16 3779 3784 3784
rect 16 13 21 3779
rect 24 3771 3776 3776
rect 24 21 29 3771
rect 32 3763 3768 3768
rect 32 29 37 3763
rect 40 3755 3760 3760
rect 40 37 45 3755
rect 48 3747 3752 3752
rect 48 45 53 3747
rect 56 3739 3744 3744
rect 56 53 61 3739
rect 64 3731 3736 3736
rect 64 61 69 3731
rect 72 3723 3728 3728
rect 72 69 77 3723
rect 80 3715 3720 3720
rect 80 77 85 3715
rect 88 3707 3712 3712
rect 88 85 93 3707
rect 96 3699 3704 3704
rect 96 93 101 3699
rect 104 3691 3696 3696
rect 104 101 109 3691
rect 112 3683 3688 3688
rect 112 109 117 3683
rect 120 3675 3680 3680
rect 120 117 125 3675
rect 128 3667 3672 3672
rect 128 125 133 3667
rect 136 3659 3664 3664
rect 136 133 141 3659
rect 144 3651 3656 3656
rect 144 141 149 3651
rect 152 3643 3648 3648
rect 152 149 157 3643
rect 160 3635 3640 3640
rect 160 157 165 3635
rect 168 3627 3632 3632
rect 168 165 173 3627
rect 176 3619 3624 3624
rect 176 173 181 3619
rect 184 3611 3616 3616
rect 184 181 189 3611
rect 192 3603 3608 3608
rect 192 189 197 3603
rect 200 3595 3600 3600
rect 200 197 205 3595
rect 208 3587 3592 3592
rect 208 205 213 3587
rect 216 3579 3584 3584
rect 216 213 221 3579
rect 224 3571 3576 3576
rect 224 221 229 3571
rect 232 3563 3568 3568
rect 232 229 237 3563
rect 240 3555 3560 3560
rect 240 237 245 3555
rect 248 3547 3552 3552
rect 248 245 253 3547
rect 256 3539 3544 3544
rect 256 253 261 3539
rect 264 3531 3536 3536
rect 264 261 269 3531
rect 272 3523 3528 3528
rect 272 269 277 3523
rect 280 3515 3520 3520
rect 280 277 285 3515
rect 288 3507 3512 3512
rect 288 285 293 3507
rect 296 3499 3504 3504
rect 296 293 301 3499
rect 304 3491 3496 3496
rect 304 301 309 3491
rect 312 3483 3488 3488
rect 312 309 317 3483
rect 320 3475 3480 3480
rect 320 317 325 3475
rect 328 3467 3472 3472
rect 328 325 333 3467
rect 336 3459 3464 3464
rect 336 333 341 3459
rect 344 3451 3456 3456
rect 344 341 349 3451
rect 352 3443 3448 3448
rect 352 349 357 3443
rect 360 3435 3440 3440
rect 360 357 365 3435
rect 368 3427 3432 3432
rect 368 365 373 3427
rect 376 3419 3424 3424
rect 376 373 381 3419
rect 384 3411 3416 3416
rect 384 381 389 3411
rect 392 3403 3408 3408
rect 392 389 397 3403
rect 400 3395 3400 3400
rect 400 397 405 3395
rect 408 3387 3392 3392
rect 408 405 413 3387
rect 416 3379 3384 3384
rect 416 413 421 3379
rect 424 3371 3376 3376
rect 424 421 429 3371
rect 432 3363 3368 3368
rect 432 429 437 3363
rect 440 3355 3360 3360
rect 440 437 445 3355
rect 448 3347 3352 3352
rect 448 445 453 3347
rect 456 3339 3344 3344
rect 456 453 461 3339
rect 464 3331 3336 3336
rect 464 461 469 3331
rect 472 3323 3328 3328
rect 472 469 477 3323
rect 480 3315 3320 3320
rect 480 477 485 3315
rect 488 3307 3312 3312
rect 488 485 493 3307
rect 496 3299 3304 3304
rect 496 493 501 3299
rect 504 3291 3296 3296
rect 504 501 509 3291
rect 512 3283 3288 3288
rect 512 509 517 3283
rect 520 3275 3280 3280
rect 520 517 525 3275
rect 528 3267 3272 3272
rect 528 525 533 3267
rect 536 3259 3264 3264
rect 536 533 541 3259
rect 544 3251 3256 3256
rect 544 541 549 3251
rect 552 3243 3248 3248
rect 552 549 557 3243
rect 560 3235 3240 3240
rect 560 557 565 3235
rect 568 3227 3232 3232
rect 568 565 573 3227
rect 576 3219 3224 3224
rect 576 573 581 3219
rect 584 3211 3216 3216
rect 584 581 589 3211
rect 592 3203 3208 3208
rect 592 589 597 3203
rect 600 3195 3200 3200
rect 600 597 605 3195
rect 608 3187 3192 3192
rect 608 605 613 3187
rect 616 3179 3184 3184
rect 616 613 621 3179
rect 624 3171 3176 3176
rect 624 621 629 3171
rect 632 3163 3168 3168
rect 632 629 637 3163
rect 640 3155 3160 3160
rect 640 637 645 3155
rect 648 3147 3152 3152
rect 648 645 653 3147
rect 656 3139 3144 3144
rect 656 653 661 3139
rect 664 3131 3136 3136
rect 664 661 669 3131
rect 672 3123 3128 3128
rect 672 669 677 3123
rect 680 3115 3120 3120
rect 680 677 685 3115
rect 688 3107 3112 3112
rect 688 685 693 3107
rect 696 3099 3104 3104
rect 696 693 701 3099
rect 704 3091 3096 3096
rect 704 701 709 3091
rect 712 3083 3088 3088
rect 712 709 717 3083
rect 720 3075 3080 3080
rect 720 717 725 3075
rect 728 3067 3072 3072
rect 728 725 733 3067
rect 736 3059 3064 3064
rect 736 733 741 3059
rect 744 3051 3056 3056
rect 744 741 749 3051
rect 752 3043 3048 3048
rect 752 749 757 3043
rect 760 3035 3040 3040
rect 760 757 765 3035
rect 768 3027 3032 3032
rect 768 765 773 3027
rect 776 3019 3024 3024
rect 776 773 781 3019
rect 784 3011 3016 3016
rect 784 781 789 3011
rect 792 3003 3008 3008
rect 792 789 797 3003
rect 800 2995 3000 3000
rect 800 797 805 2995
rect 808 2987 2992 2992
rect 808 805 813 2987
rect 816 2979 2984 2984
rect 816 813 821 2979
rect 824 2971 2976 2976
rect 824 821 829 2971
rect 832 2963 2968 2968
rect 832 829 837 2963
rect 840 2955 2960 2960
rect 840 837 845 2955
rect 848 2947 2952 2952
rect 848 845 853 2947
rect 856 2939 2944 2944
rect 856 853 861 2939
rect 864 2931 2936 2936
rect 864 861 869 2931
rect 872 2923 2928 2928
rect 872 869 877 2923
rect 880 2915 2920 2920
rect 880 877 885 2915
rect 888 2907 2912 2912
rect 888 885 893 2907
rect 896 2899 2904 2904
rect 896 893 901 2899
rect 904 2891 2896 2896
rect 904 901 909 2891
rect 912 2883 2888 2888
rect 912 909 917 2883
rect 920 2875 2880 2880
rect 920 917 925 2875
rect 928 2867 2872 2872
rect 928 925 933 2867
rect 936 2859 2864 2864
rect 936 933 941 2859
rect 944 2851 2856 2856
rect 944 941 949 2851
rect 952 2843 2848 2848
rect 952 949 957 2843
rect 960 2835 2840 2840
rect 960 957 965 2835
rect 968 2827 2832 2832
rect 968 965 973 2827
rect 976 2819 2824 2824
rect 976 973 981 2819
rect 984 2811 2816 2816
rect 984 981 989 2811
rect 992 2803 2808 2808
rect 992 989 997 2803
rect 1000 2795 2800 2800
rect 1000 997 1005 2795
rect 1008 2787 2792 2792
rect 1008 1005 1013 2787
rect 1016 2779 2784 2784
rect 1016 1013 1021 2779
rect 1024 2771 2776 2776
rect 1024 1021 1029 2771
rect 1032 2763 2768 2768
rect 1032 1029 1037 2763
rect 1040 2755 2760 2760
rect 1040 1037 1045 2755
rect 1048 2747 2752 2752
rect 1048 1045 1053 2747
rect 1056 2739 2744 2744
rect 1056 1053 1061 2739
rect 1064 2731 2736 2736
rect 1064 1061 1069 2731
rect 1072 2723 2728 2728
rect 1072 1069 1077 2723
rect 1080 2715 2720 2720
rect 1080 1077 1085 2715
rect 1088 2707 2712 2712
rect 1088 1085 1093 2707
rect 1096 2699 2704 2704
rect 1096 1093 1101 2699
rect 1104 2691 2696 2696
rect 1104 1101 1109 2691
rect 1112 2683 2688 2688
rect 1112 1109 1117 2683
rect 1120 2675 2680 2680
rect 1120 1117 1125 2675
rect 1128 2667 2672 2672
rect 1128 1125 1133 2667
rect 1136 2659 2664 2664
rect 1136 1133 1141 2659
rect 1144 2651 2656 2656
rect 1144 1141 1149 2651
rect 1152 2643 2648 2648
rect 1152 1149 1157 2643
rect 1160 2635 2640 2640
rect 1160 1157 1165 2635
rect 1168 2627 2632 2632
rect 1168 1165 1173 2627
rect 1176 2619 2624 2624
rect 1176 1173 1181 2619
rect 1184 2611 2616 2616
rect 1184 1181 1189 2611
rect 1192 2603 2608 2608
rect 1192 1189 1197 2603
rect 1200 2595 2600 2600
rect 1200 1197 1205 2595
rect 1208 2587 2592 2592
rect 1208 1205 1213 2587
rect 1216 2579 2584 2584
rect 1216 1213 1221 2579
rect 1224 2571 2576 2576
rect 1224 1221 1229 2571
rect 1232 2563 2568 2568
rect 1232 1229 1237 2563
rect 1240 2555 2560 2560
rect 1240 1237 1245 2555
rect 1248 2547 2552 2552
rect 1248 1245 1253 2547
rect 1256 2539 2544 2544
rect 1256 1253 1261 2539
rect 1264 2531 2536 2536
rect 1264 1261 1269 2531
rect 1272 2523 2528 2528
rect 1272 1269 1277 2523
rect 1280 2515 2520 2520
rect 1280 1277 1285 2515
rect 1288 2507 2512 2512
rect 1288 1285 1293 2507
rect 1296 2499 2504 2504
rect 1296 1293 1301 2499
rect 1304 2491 2496 2496
rect 1304 1301 1309 2491
rect 1312 2483 2488 2488
rect 1312 1309 1317 2483
rect 1320 2475 2480 2480
rect 1320 1317 1325 2475
rect 1328 2467 2472 2472
rect 1328 1325 1333 2467
rect 1336 2459 2464 2464
rect 1336 1333 1341 2459
rect 1344 2451 2456 2456
rect 1344 1341 1349 2451
rect 1352 2443 2448 2448
rect 1352 1349 1357 2443
rect 1360 2435 2440 2440
rect 1360 1357 1365 2435
rect 1368 2427 2432 2432
rect 1368 1365 1373 2427
rect 1376 2419 2424 2424
rect 1376 1373 1381 2419
rect 1384 2411 2416 2416
rect 1384 1381 1389 2411
rect 1392 2403 2408 2408
rect 1392 1389 1397 2403
rect 1400 2395 2400 2400
rect 1400 1397 1405 2395
rect 1408 2387 2392 2392
rect 1408 1405 1413 2387
rect 1416 2379 2384 2384
rect 1416 1413 1421 2379
rect 1424 2371 2376 2376
rect 1424 1421 1429 2371
rect 1432 2363 2368 2368
rect 1432 1429 1437 2363
rect 1440 2355 2360 2360
rect 1440 1437 1445 2355
rect 1448 2347 2352 2352
rect 1448 1445 1453 2347
rect 1456 2339 2344 2344
rect 1456 1453 1461 2339
rect 1464 2331 2336 2336
rect 1464 1461 1469 2331
rect 1472 2323 2328 2328
rect 1472 1469 1477 2323
rect 1480 2315 2320 2320
rect 1480 1477 1485 2315
rect 1488 2307 2312 2312
rect 1488 1485 1493 2307
rect 1496 2299 2304 2304
rect 1496 1493 1501 2299
rect 1504 2291 2296 2296
rect 1504 1501 1509 2291
rect 1512 2283 2288 2288
rect 1512 1509 1517 2283
rect 1520 2275 2280 2280
rect 1520 1517 1525 2275
rect 1528 2267 2272 2272
rect 1528 1525 1533 2267
rect 1536 2259 2264 2264
rect 1536 1533 1541 2259
rect 1544 2251 2256 2256
rect 1544 1541 1549 2251
rect 1552 2243 2248 2248
rect 1552 1549 1557 2243
rect 1560 2235 2240 2240
rect 1560 1557 1565 2235
rect 1568 2227 2232 2232
rect 1568 1565 1573 2227
rect 1576 2219 2224 2224
rect 1576 1573 1581 2219
rect 1584 2211 2216 2216
rect 1584 1581 1589 2211
rect 1592 2203 2208 2208
rect 1592 1589 1597 2203
rect 1600 2195 2200 2200
rect 1600 1597 1605 2195
rect 1608 2187 2192 2192
rect 1608 1605 1613 2187
rect 1616 2179 2184 2184
rect 1616 1613 1621 2179
rect 1624 2171 2176 2176
rect 1624 1621 1629 2171
rect 1632 2163 2168 2168
rect 1632 1629 1637 2163
rect 1640 2155 2160 2160
rect 1640 1637 1645 2155
rect 1648 2147 2152 2152
rect 1648 1645 1653 2147
rect 1656 2139 2144 2144
rect 1656 1653 1661 2139
rect 1664 2131 2136 2136
rect 1664 1661 1669 2131
rect 1672 2123 2128 2128
rect 1672 1669 1677 2123
rect 1680 2115 2120 2120
rect 1680 1677 1685 2115
rect 1688 2107 2112 2112
rect 1688 1685 1693 2107
rect 1696 2099 2104 2104
rect 1696 1693 1701 2099
rect 1704 2091 2096 2096
rect 1704 1701 1709 2091
rect 1712 2083 2088 2088
rect 1712 1709 1717 2083
rect 1720 2075 2080 2080
rect 1720 1717 1725 2075
rect 1728 2067 2072 2072
rect 1728 1725 1733 2067
rect 1736 2059 2064 2064
rect 1736 1733 1741 2059
rect 1744 2051 2056 2056
rect 1744 1741 1749 2051
rect 1752 2043 2048 2048
rect 1752 1749 1757 2043
rect 1760 2035 2040 2040
rect 1760 1757 1765 2035
rect 1768 2027 2032 2032
rect 1768 1765 1773 2027
rect 1776 2019 2024 2024
rect 1776 1773 1781 2019
rect 1784 2011 2016 2016
rect 1784 1781 1789 2011
rect 1792 2003 2008 2008
rect 1792 1789 1797 2003
rect 1800 1995 2000 2000
rect 1800 1797 1805 1995
rect 1808 1987 1992 1992
rect 1808 1805 1813 1987
rect 1816 1979 1984 1984
rect 1816 1813 1821 1979
rect 1824 1971 1976 1976
rect 1824 1821 1829 1971
rect 1832 1963 1968 1968
rect 1832 1829 1837 1963
rect 1840 1955 1960 1960
rect 1840 1837 1845 1955
rect 1848 1947 1952 1952
rect 1848 1845 1853 1947
rect 1856 1939 1944 1944
rect 1856 1853 1861 1939
rect 1864 1931 1936 1936
rect 1864 1861 1869 1931
rect 1872 1923 1928 1928
rect 1872 1869 1877 1923
rect 1880 1915 1920 1920
rect 1880 1877 1885 1915
rect 1888 1907 1912 1912
rect 1888 1885 1893 1907
rect 1896 1894 1903 1895
rect 1896 1889 1897 1894
rect 1902 1893 1903 1894
rect 1907 1893 1912 1907
rect 1902 1889 1912 1893
rect 1896 1888 1912 1889
rect 1915 1885 1920 1915
rect 1888 1880 1920 1885
rect 1923 1877 1928 1923
rect 1880 1872 1928 1877
rect 1931 1869 1936 1931
rect 1872 1864 1936 1869
rect 1939 1861 1944 1939
rect 1864 1856 1944 1861
rect 1947 1853 1952 1947
rect 1856 1848 1952 1853
rect 1955 1845 1960 1955
rect 1848 1840 1960 1845
rect 1963 1837 1968 1963
rect 1840 1832 1968 1837
rect 1971 1829 1976 1971
rect 1832 1824 1976 1829
rect 1979 1821 1984 1979
rect 1824 1816 1984 1821
rect 1987 1813 1992 1987
rect 1816 1808 1992 1813
rect 1995 1805 2000 1995
rect 1808 1800 2000 1805
rect 2003 1797 2008 2003
rect 1800 1792 2008 1797
rect 2011 1789 2016 2011
rect 1792 1784 2016 1789
rect 2019 1781 2024 2019
rect 1784 1776 2024 1781
rect 2027 1773 2032 2027
rect 1776 1768 2032 1773
rect 2035 1765 2040 2035
rect 1768 1760 2040 1765
rect 2043 1757 2048 2043
rect 1760 1752 2048 1757
rect 2051 1749 2056 2051
rect 1752 1744 2056 1749
rect 2059 1741 2064 2059
rect 1744 1736 2064 1741
rect 2067 1733 2072 2067
rect 1736 1728 2072 1733
rect 2075 1725 2080 2075
rect 1728 1720 2080 1725
rect 2083 1717 2088 2083
rect 1720 1712 2088 1717
rect 2091 1709 2096 2091
rect 1712 1704 2096 1709
rect 2099 1701 2104 2099
rect 1704 1696 2104 1701
rect 2107 1693 2112 2107
rect 1696 1688 2112 1693
rect 2115 1685 2120 2115
rect 1688 1680 2120 1685
rect 2123 1677 2128 2123
rect 1680 1672 2128 1677
rect 2131 1669 2136 2131
rect 1672 1664 2136 1669
rect 2139 1661 2144 2139
rect 1664 1656 2144 1661
rect 2147 1653 2152 2147
rect 1656 1648 2152 1653
rect 2155 1645 2160 2155
rect 1648 1640 2160 1645
rect 2163 1637 2168 2163
rect 1640 1632 2168 1637
rect 2171 1629 2176 2171
rect 1632 1624 2176 1629
rect 2179 1621 2184 2179
rect 1624 1616 2184 1621
rect 2187 1613 2192 2187
rect 1616 1608 2192 1613
rect 2195 1605 2200 2195
rect 1608 1600 2200 1605
rect 2203 1597 2208 2203
rect 1600 1592 2208 1597
rect 2211 1589 2216 2211
rect 1592 1584 2216 1589
rect 2219 1581 2224 2219
rect 1584 1576 2224 1581
rect 2227 1573 2232 2227
rect 1576 1568 2232 1573
rect 2235 1565 2240 2235
rect 1568 1560 2240 1565
rect 2243 1557 2248 2243
rect 1560 1552 2248 1557
rect 2251 1549 2256 2251
rect 1552 1544 2256 1549
rect 2259 1541 2264 2259
rect 1544 1536 2264 1541
rect 2267 1533 2272 2267
rect 1536 1528 2272 1533
rect 2275 1525 2280 2275
rect 1528 1520 2280 1525
rect 2283 1517 2288 2283
rect 1520 1512 2288 1517
rect 2291 1509 2296 2291
rect 1512 1504 2296 1509
rect 2299 1501 2304 2299
rect 1504 1496 2304 1501
rect 2307 1493 2312 2307
rect 1496 1488 2312 1493
rect 2315 1485 2320 2315
rect 1488 1480 2320 1485
rect 2323 1477 2328 2323
rect 1480 1472 2328 1477
rect 2331 1469 2336 2331
rect 1472 1464 2336 1469
rect 2339 1461 2344 2339
rect 1464 1456 2344 1461
rect 2347 1453 2352 2347
rect 1456 1448 2352 1453
rect 2355 1445 2360 2355
rect 1448 1440 2360 1445
rect 2363 1437 2368 2363
rect 1440 1432 2368 1437
rect 2371 1429 2376 2371
rect 1432 1424 2376 1429
rect 2379 1421 2384 2379
rect 1424 1416 2384 1421
rect 2387 1413 2392 2387
rect 1416 1408 2392 1413
rect 2395 1405 2400 2395
rect 1408 1400 2400 1405
rect 2403 1397 2408 2403
rect 1400 1392 2408 1397
rect 2411 1389 2416 2411
rect 1392 1384 2416 1389
rect 2419 1381 2424 2419
rect 1384 1376 2424 1381
rect 2427 1373 2432 2427
rect 1376 1368 2432 1373
rect 2435 1365 2440 2435
rect 1368 1360 2440 1365
rect 2443 1357 2448 2443
rect 1360 1352 2448 1357
rect 2451 1349 2456 2451
rect 1352 1344 2456 1349
rect 2459 1341 2464 2459
rect 1344 1336 2464 1341
rect 2467 1333 2472 2467
rect 1336 1328 2472 1333
rect 2475 1325 2480 2475
rect 1328 1320 2480 1325
rect 2483 1317 2488 2483
rect 1320 1312 2488 1317
rect 2491 1309 2496 2491
rect 1312 1304 2496 1309
rect 2499 1301 2504 2499
rect 1304 1296 2504 1301
rect 2507 1293 2512 2507
rect 1296 1288 2512 1293
rect 2515 1285 2520 2515
rect 1288 1280 2520 1285
rect 2523 1277 2528 2523
rect 1280 1272 2528 1277
rect 2531 1269 2536 2531
rect 1272 1264 2536 1269
rect 2539 1261 2544 2539
rect 1264 1256 2544 1261
rect 2547 1253 2552 2547
rect 1256 1248 2552 1253
rect 2555 1245 2560 2555
rect 1248 1240 2560 1245
rect 2563 1237 2568 2563
rect 1240 1232 2568 1237
rect 2571 1229 2576 2571
rect 1232 1224 2576 1229
rect 2579 1221 2584 2579
rect 1224 1216 2584 1221
rect 2587 1213 2592 2587
rect 1216 1208 2592 1213
rect 2595 1205 2600 2595
rect 1208 1200 2600 1205
rect 2603 1197 2608 2603
rect 1200 1192 2608 1197
rect 2611 1189 2616 2611
rect 1192 1184 2616 1189
rect 2619 1181 2624 2619
rect 1184 1176 2624 1181
rect 2627 1173 2632 2627
rect 1176 1168 2632 1173
rect 2635 1165 2640 2635
rect 1168 1160 2640 1165
rect 2643 1157 2648 2643
rect 1160 1152 2648 1157
rect 2651 1149 2656 2651
rect 1152 1144 2656 1149
rect 2659 1141 2664 2659
rect 1144 1136 2664 1141
rect 2667 1133 2672 2667
rect 1136 1128 2672 1133
rect 2675 1125 2680 2675
rect 1128 1120 2680 1125
rect 2683 1117 2688 2683
rect 1120 1112 2688 1117
rect 2691 1109 2696 2691
rect 1112 1104 2696 1109
rect 2699 1101 2704 2699
rect 1104 1096 2704 1101
rect 2707 1093 2712 2707
rect 1096 1088 2712 1093
rect 2715 1085 2720 2715
rect 1088 1080 2720 1085
rect 2723 1077 2728 2723
rect 1080 1072 2728 1077
rect 2731 1069 2736 2731
rect 1072 1064 2736 1069
rect 2739 1061 2744 2739
rect 1064 1056 2744 1061
rect 2747 1053 2752 2747
rect 1056 1048 2752 1053
rect 2755 1045 2760 2755
rect 1048 1040 2760 1045
rect 2763 1037 2768 2763
rect 1040 1032 2768 1037
rect 2771 1029 2776 2771
rect 1032 1024 2776 1029
rect 2779 1021 2784 2779
rect 1024 1016 2784 1021
rect 2787 1013 2792 2787
rect 1016 1008 2792 1013
rect 2795 1005 2800 2795
rect 1008 1000 2800 1005
rect 2803 997 2808 2803
rect 1000 992 2808 997
rect 2811 989 2816 2811
rect 992 984 2816 989
rect 2819 981 2824 2819
rect 984 976 2824 981
rect 2827 973 2832 2827
rect 976 968 2832 973
rect 2835 965 2840 2835
rect 968 960 2840 965
rect 2843 957 2848 2843
rect 960 952 2848 957
rect 2851 949 2856 2851
rect 952 944 2856 949
rect 2859 941 2864 2859
rect 944 936 2864 941
rect 2867 933 2872 2867
rect 936 928 2872 933
rect 2875 925 2880 2875
rect 928 920 2880 925
rect 2883 917 2888 2883
rect 920 912 2888 917
rect 2891 909 2896 2891
rect 912 904 2896 909
rect 2899 901 2904 2899
rect 904 896 2904 901
rect 2907 893 2912 2907
rect 896 888 2912 893
rect 2915 885 2920 2915
rect 888 880 2920 885
rect 2923 877 2928 2923
rect 880 872 2928 877
rect 2931 869 2936 2931
rect 872 864 2936 869
rect 2939 861 2944 2939
rect 864 856 2944 861
rect 2947 853 2952 2947
rect 856 848 2952 853
rect 2955 845 2960 2955
rect 848 840 2960 845
rect 2963 837 2968 2963
rect 840 832 2968 837
rect 2971 829 2976 2971
rect 832 824 2976 829
rect 2979 821 2984 2979
rect 824 816 2984 821
rect 2987 813 2992 2987
rect 816 808 2992 813
rect 2995 805 3000 2995
rect 808 800 3000 805
rect 3003 797 3008 3003
rect 800 792 3008 797
rect 3011 789 3016 3011
rect 792 784 3016 789
rect 3019 781 3024 3019
rect 784 776 3024 781
rect 3027 773 3032 3027
rect 776 768 3032 773
rect 3035 765 3040 3035
rect 768 760 3040 765
rect 3043 757 3048 3043
rect 760 752 3048 757
rect 3051 749 3056 3051
rect 752 744 3056 749
rect 3059 741 3064 3059
rect 744 736 3064 741
rect 3067 733 3072 3067
rect 736 728 3072 733
rect 3075 725 3080 3075
rect 728 720 3080 725
rect 3083 717 3088 3083
rect 720 712 3088 717
rect 3091 709 3096 3091
rect 712 704 3096 709
rect 3099 701 3104 3099
rect 704 696 3104 701
rect 3107 693 3112 3107
rect 696 688 3112 693
rect 3115 685 3120 3115
rect 688 680 3120 685
rect 3123 677 3128 3123
rect 680 672 3128 677
rect 3131 669 3136 3131
rect 672 664 3136 669
rect 3139 661 3144 3139
rect 664 656 3144 661
rect 3147 653 3152 3147
rect 656 648 3152 653
rect 3155 645 3160 3155
rect 648 640 3160 645
rect 3163 637 3168 3163
rect 640 632 3168 637
rect 3171 629 3176 3171
rect 632 624 3176 629
rect 3179 621 3184 3179
rect 624 616 3184 621
rect 3187 613 3192 3187
rect 616 608 3192 613
rect 3195 605 3200 3195
rect 608 600 3200 605
rect 3203 597 3208 3203
rect 600 592 3208 597
rect 3211 589 3216 3211
rect 592 584 3216 589
rect 3219 581 3224 3219
rect 584 576 3224 581
rect 3227 573 3232 3227
rect 576 568 3232 573
rect 3235 565 3240 3235
rect 568 560 3240 565
rect 3243 557 3248 3243
rect 560 552 3248 557
rect 3251 549 3256 3251
rect 552 544 3256 549
rect 3259 541 3264 3259
rect 544 536 3264 541
rect 3267 533 3272 3267
rect 536 528 3272 533
rect 3275 525 3280 3275
rect 528 520 3280 525
rect 3283 517 3288 3283
rect 520 512 3288 517
rect 3291 509 3296 3291
rect 512 504 3296 509
rect 3299 501 3304 3299
rect 504 496 3304 501
rect 3307 493 3312 3307
rect 496 488 3312 493
rect 3315 485 3320 3315
rect 488 480 3320 485
rect 3323 477 3328 3323
rect 480 472 3328 477
rect 3331 469 3336 3331
rect 472 464 3336 469
rect 3339 461 3344 3339
rect 464 456 3344 461
rect 3347 453 3352 3347
rect 456 448 3352 453
rect 3355 445 3360 3355
rect 448 440 3360 445
rect 3363 437 3368 3363
rect 440 432 3368 437
rect 3371 429 3376 3371
rect 432 424 3376 429
rect 3379 421 3384 3379
rect 424 416 3384 421
rect 3387 413 3392 3387
rect 416 408 3392 413
rect 3395 405 3400 3395
rect 408 400 3400 405
rect 3403 397 3408 3403
rect 400 392 3408 397
rect 3411 389 3416 3411
rect 392 384 3416 389
rect 3419 381 3424 3419
rect 384 376 3424 381
rect 3427 373 3432 3427
rect 376 368 3432 373
rect 3435 365 3440 3435
rect 368 360 3440 365
rect 3443 357 3448 3443
rect 360 352 3448 357
rect 3451 349 3456 3451
rect 352 344 3456 349
rect 3459 341 3464 3459
rect 344 336 3464 341
rect 3467 333 3472 3467
rect 336 328 3472 333
rect 3475 325 3480 3475
rect 328 320 3480 325
rect 3483 317 3488 3483
rect 320 312 3488 317
rect 3491 309 3496 3491
rect 312 304 3496 309
rect 3499 301 3504 3499
rect 304 296 3504 301
rect 3507 293 3512 3507
rect 296 288 3512 293
rect 3515 285 3520 3515
rect 288 280 3520 285
rect 3523 277 3528 3523
rect 280 272 3528 277
rect 3531 269 3536 3531
rect 272 264 3536 269
rect 3539 261 3544 3539
rect 264 256 3544 261
rect 3547 253 3552 3547
rect 256 248 3552 253
rect 3555 245 3560 3555
rect 248 240 3560 245
rect 3563 237 3568 3563
rect 240 232 3568 237
rect 3571 229 3576 3571
rect 232 224 3576 229
rect 3579 221 3584 3579
rect 224 216 3584 221
rect 3587 213 3592 3587
rect 216 208 3592 213
rect 3595 205 3600 3595
rect 208 200 3600 205
rect 3603 197 3608 3603
rect 200 192 3608 197
rect 3611 189 3616 3611
rect 192 184 3616 189
rect 3619 181 3624 3619
rect 184 176 3624 181
rect 3627 173 3632 3627
rect 176 168 3632 173
rect 3635 165 3640 3635
rect 168 160 3640 165
rect 3643 157 3648 3643
rect 160 152 3648 157
rect 3651 149 3656 3651
rect 152 144 3656 149
rect 3659 141 3664 3659
rect 144 136 3664 141
rect 3667 133 3672 3667
rect 136 128 3672 133
rect 3675 125 3680 3675
rect 128 120 3680 125
rect 3683 117 3688 3683
rect 120 112 3688 117
rect 3691 109 3696 3691
rect 112 104 3696 109
rect 3699 101 3704 3699
rect 104 96 3704 101
rect 3707 93 3712 3707
rect 96 88 3712 93
rect 3715 85 3720 3715
rect 88 80 3720 85
rect 3723 77 3728 3723
rect 80 72 3728 77
rect 3731 69 3736 3731
rect 72 64 3736 69
rect 3739 61 3744 3739
rect 64 56 3744 61
rect 3747 53 3752 3747
rect 56 48 3752 53
rect 3755 45 3760 3755
rect 48 40 3760 45
rect 3763 37 3768 3763
rect 40 32 3768 37
rect 3771 29 3776 3771
rect 32 24 3776 29
rect 3779 21 3784 3779
rect 24 16 3784 21
rect 3787 13 3792 3787
rect 16 8 3792 13
rect 3795 5 3800 3795
rect 8 0 3800 5
rect -1 -1 5 0
<< end >>
