magic
tech scmos
timestamp 1417795444
<< nwell >>
rect 150 -149 300 -75
<< ntransistor >>
rect 163 -162 165 -156
rect 171 -162 173 -156
rect 179 -162 181 -156
rect 197 -186 199 -156
rect 214 -186 216 -156
rect 222 -186 224 -156
rect 230 -186 232 -156
rect 238 -186 240 -156
rect 246 -186 248 -156
rect 254 -186 256 -156
rect 262 -186 264 -156
rect 270 -186 272 -156
rect 278 -186 280 -156
rect 286 -186 288 -156
<< ptransistor >>
rect 163 -141 165 -135
rect 168 -141 170 -135
rect 177 -141 179 -135
rect 197 -141 199 -81
rect 214 -141 216 -81
rect 222 -141 224 -81
rect 230 -141 232 -81
rect 238 -141 240 -81
rect 246 -141 248 -81
rect 254 -141 256 -81
rect 262 -141 264 -81
rect 270 -141 272 -81
rect 278 -141 280 -81
rect 286 -141 288 -81
<< ndiffusion >>
rect 157 -157 163 -156
rect 157 -161 158 -157
rect 162 -161 163 -157
rect 157 -162 163 -161
rect 165 -157 171 -156
rect 165 -161 166 -157
rect 170 -161 171 -157
rect 165 -162 171 -161
rect 173 -157 179 -156
rect 173 -161 174 -157
rect 178 -161 179 -157
rect 173 -162 179 -161
rect 181 -157 187 -156
rect 181 -161 182 -157
rect 186 -161 187 -157
rect 181 -162 187 -161
rect 191 -157 197 -156
rect 191 -161 192 -157
rect 196 -161 197 -157
rect 191 -165 197 -161
rect 191 -169 192 -165
rect 196 -169 197 -165
rect 191 -173 197 -169
rect 191 -177 192 -173
rect 196 -177 197 -173
rect 191 -181 197 -177
rect 191 -185 192 -181
rect 196 -185 197 -181
rect 191 -186 197 -185
rect 199 -157 205 -156
rect 199 -185 200 -157
rect 204 -185 205 -157
rect 199 -186 205 -185
rect 208 -157 214 -156
rect 208 -161 209 -157
rect 213 -161 214 -157
rect 208 -165 214 -161
rect 208 -169 209 -165
rect 213 -169 214 -165
rect 208 -173 214 -169
rect 208 -177 209 -173
rect 213 -177 214 -173
rect 208 -181 214 -177
rect 208 -185 209 -181
rect 213 -185 214 -181
rect 208 -186 214 -185
rect 216 -157 222 -156
rect 216 -185 217 -157
rect 221 -185 222 -157
rect 216 -186 222 -185
rect 224 -157 230 -156
rect 224 -161 225 -157
rect 229 -161 230 -157
rect 224 -165 230 -161
rect 224 -169 225 -165
rect 229 -169 230 -165
rect 224 -173 230 -169
rect 224 -177 225 -173
rect 229 -177 230 -173
rect 224 -181 230 -177
rect 224 -185 225 -181
rect 229 -185 230 -181
rect 224 -186 230 -185
rect 232 -157 238 -156
rect 232 -185 233 -157
rect 237 -185 238 -157
rect 232 -186 238 -185
rect 240 -157 246 -156
rect 240 -161 241 -157
rect 245 -161 246 -157
rect 240 -165 246 -161
rect 240 -169 241 -165
rect 245 -169 246 -165
rect 240 -173 246 -169
rect 240 -177 241 -173
rect 245 -177 246 -173
rect 240 -181 246 -177
rect 240 -185 241 -181
rect 245 -185 246 -181
rect 240 -186 246 -185
rect 248 -157 254 -156
rect 248 -185 249 -157
rect 253 -185 254 -157
rect 248 -186 254 -185
rect 256 -157 262 -156
rect 256 -161 257 -157
rect 261 -161 262 -157
rect 256 -165 262 -161
rect 256 -169 257 -165
rect 261 -169 262 -165
rect 256 -173 262 -169
rect 256 -177 257 -173
rect 261 -177 262 -173
rect 256 -181 262 -177
rect 256 -185 257 -181
rect 261 -185 262 -181
rect 256 -186 262 -185
rect 264 -157 270 -156
rect 264 -185 265 -157
rect 269 -185 270 -157
rect 264 -186 270 -185
rect 272 -157 278 -156
rect 272 -161 273 -157
rect 277 -161 278 -157
rect 272 -165 278 -161
rect 272 -169 273 -165
rect 277 -169 278 -165
rect 272 -173 278 -169
rect 272 -177 273 -173
rect 277 -177 278 -173
rect 272 -181 278 -177
rect 272 -185 273 -181
rect 277 -185 278 -181
rect 272 -186 278 -185
rect 280 -157 286 -156
rect 280 -185 281 -157
rect 285 -185 286 -157
rect 280 -186 286 -185
rect 288 -157 294 -156
rect 288 -161 289 -157
rect 293 -161 294 -157
rect 288 -165 294 -161
rect 288 -169 289 -165
rect 293 -169 294 -165
rect 288 -173 294 -169
rect 288 -177 289 -173
rect 293 -177 294 -173
rect 288 -181 294 -177
rect 288 -185 289 -181
rect 293 -185 294 -181
rect 288 -186 294 -185
<< pdiffusion >>
rect 191 -82 197 -81
rect 191 -86 192 -82
rect 196 -86 197 -82
rect 191 -90 197 -86
rect 191 -94 192 -90
rect 196 -94 197 -90
rect 191 -98 197 -94
rect 191 -102 192 -98
rect 196 -102 197 -98
rect 191 -106 197 -102
rect 191 -116 192 -106
rect 196 -116 197 -106
rect 191 -120 197 -116
rect 191 -124 192 -120
rect 196 -124 197 -120
rect 191 -128 197 -124
rect 191 -132 192 -128
rect 196 -132 197 -128
rect 157 -136 163 -135
rect 157 -140 158 -136
rect 162 -140 163 -136
rect 157 -141 163 -140
rect 165 -141 168 -135
rect 170 -136 177 -135
rect 170 -140 171 -136
rect 175 -140 177 -136
rect 170 -141 177 -140
rect 179 -136 185 -135
rect 179 -140 180 -136
rect 184 -140 185 -136
rect 179 -141 185 -140
rect 191 -136 197 -132
rect 191 -140 192 -136
rect 196 -140 197 -136
rect 191 -141 197 -140
rect 199 -82 205 -81
rect 199 -140 200 -82
rect 204 -140 205 -82
rect 199 -141 205 -140
rect 208 -82 214 -81
rect 208 -86 209 -82
rect 213 -86 214 -82
rect 208 -90 214 -86
rect 208 -94 209 -90
rect 213 -94 214 -90
rect 208 -98 214 -94
rect 208 -102 209 -98
rect 213 -102 214 -98
rect 208 -106 214 -102
rect 208 -116 209 -106
rect 213 -116 214 -106
rect 208 -120 214 -116
rect 208 -124 209 -120
rect 213 -124 214 -120
rect 208 -128 214 -124
rect 208 -132 209 -128
rect 213 -132 214 -128
rect 208 -136 214 -132
rect 208 -140 209 -136
rect 213 -140 214 -136
rect 208 -141 214 -140
rect 216 -82 222 -81
rect 216 -140 217 -82
rect 221 -140 222 -82
rect 216 -141 222 -140
rect 224 -82 230 -81
rect 224 -86 225 -82
rect 229 -86 230 -82
rect 224 -90 230 -86
rect 224 -94 225 -90
rect 229 -94 230 -90
rect 224 -98 230 -94
rect 224 -102 225 -98
rect 229 -102 230 -98
rect 224 -106 230 -102
rect 224 -116 225 -106
rect 229 -116 230 -106
rect 224 -120 230 -116
rect 224 -124 225 -120
rect 229 -124 230 -120
rect 224 -128 230 -124
rect 224 -132 225 -128
rect 229 -132 230 -128
rect 224 -136 230 -132
rect 224 -140 225 -136
rect 229 -140 230 -136
rect 224 -141 230 -140
rect 232 -82 238 -81
rect 232 -140 233 -82
rect 237 -140 238 -82
rect 232 -141 238 -140
rect 240 -82 246 -81
rect 240 -86 241 -82
rect 245 -86 246 -82
rect 240 -90 246 -86
rect 240 -94 241 -90
rect 245 -94 246 -90
rect 240 -98 246 -94
rect 240 -102 241 -98
rect 245 -102 246 -98
rect 240 -106 246 -102
rect 240 -116 241 -106
rect 245 -116 246 -106
rect 240 -120 246 -116
rect 240 -124 241 -120
rect 245 -124 246 -120
rect 240 -128 246 -124
rect 240 -132 241 -128
rect 245 -132 246 -128
rect 240 -136 246 -132
rect 240 -140 241 -136
rect 245 -140 246 -136
rect 240 -141 246 -140
rect 248 -82 254 -81
rect 248 -140 249 -82
rect 253 -140 254 -82
rect 248 -141 254 -140
rect 256 -82 262 -81
rect 256 -86 257 -82
rect 261 -86 262 -82
rect 256 -90 262 -86
rect 256 -94 257 -90
rect 261 -94 262 -90
rect 256 -98 262 -94
rect 256 -102 257 -98
rect 261 -102 262 -98
rect 256 -106 262 -102
rect 256 -116 257 -106
rect 261 -116 262 -106
rect 256 -120 262 -116
rect 256 -124 257 -120
rect 261 -124 262 -120
rect 256 -128 262 -124
rect 256 -132 257 -128
rect 261 -132 262 -128
rect 256 -136 262 -132
rect 256 -140 257 -136
rect 261 -140 262 -136
rect 256 -141 262 -140
rect 264 -82 270 -81
rect 264 -140 265 -82
rect 269 -140 270 -82
rect 264 -141 270 -140
rect 272 -82 278 -81
rect 272 -86 273 -82
rect 277 -86 278 -82
rect 272 -90 278 -86
rect 272 -94 273 -90
rect 277 -94 278 -90
rect 272 -98 278 -94
rect 272 -102 273 -98
rect 277 -102 278 -98
rect 272 -106 278 -102
rect 272 -116 273 -106
rect 277 -116 278 -106
rect 272 -120 278 -116
rect 272 -124 273 -120
rect 277 -124 278 -120
rect 272 -128 278 -124
rect 272 -132 273 -128
rect 277 -132 278 -128
rect 272 -136 278 -132
rect 272 -140 273 -136
rect 277 -140 278 -136
rect 272 -141 278 -140
rect 280 -82 286 -81
rect 280 -140 281 -82
rect 285 -140 286 -82
rect 280 -141 286 -140
rect 288 -82 294 -81
rect 288 -86 289 -82
rect 293 -86 294 -82
rect 288 -90 294 -86
rect 288 -94 289 -90
rect 293 -94 294 -90
rect 288 -98 294 -94
rect 288 -102 289 -98
rect 293 -102 294 -98
rect 288 -106 294 -102
rect 288 -116 289 -106
rect 293 -116 294 -106
rect 288 -120 294 -116
rect 288 -124 289 -120
rect 293 -124 294 -120
rect 288 -128 294 -124
rect 288 -132 289 -128
rect 293 -132 294 -128
rect 288 -136 294 -132
rect 288 -140 289 -136
rect 293 -140 294 -136
rect 288 -141 294 -140
<< ndcontact >>
rect 158 -161 162 -157
rect 166 -161 170 -157
rect 174 -161 178 -157
rect 182 -161 186 -157
rect 192 -161 196 -157
rect 192 -169 196 -165
rect 192 -177 196 -173
rect 192 -185 196 -181
rect 200 -185 204 -157
rect 209 -161 213 -157
rect 209 -169 213 -165
rect 209 -177 213 -173
rect 209 -185 213 -181
rect 217 -185 221 -157
rect 225 -161 229 -157
rect 225 -169 229 -165
rect 225 -177 229 -173
rect 225 -185 229 -181
rect 233 -185 237 -157
rect 241 -161 245 -157
rect 241 -169 245 -165
rect 241 -177 245 -173
rect 241 -185 245 -181
rect 249 -185 253 -157
rect 257 -161 261 -157
rect 257 -169 261 -165
rect 257 -177 261 -173
rect 257 -185 261 -181
rect 265 -185 269 -157
rect 273 -161 277 -157
rect 273 -169 277 -165
rect 273 -177 277 -173
rect 273 -185 277 -181
rect 281 -185 285 -157
rect 289 -161 293 -157
rect 289 -169 293 -165
rect 289 -177 293 -173
rect 289 -185 293 -181
<< pdcontact >>
rect 192 -86 196 -82
rect 192 -94 196 -90
rect 192 -102 196 -98
rect 192 -116 196 -106
rect 192 -124 196 -120
rect 192 -132 196 -128
rect 158 -140 162 -136
rect 171 -140 175 -136
rect 180 -140 184 -136
rect 192 -140 196 -136
rect 200 -140 204 -82
rect 209 -86 213 -82
rect 209 -94 213 -90
rect 209 -102 213 -98
rect 209 -116 213 -106
rect 209 -124 213 -120
rect 209 -132 213 -128
rect 209 -140 213 -136
rect 217 -140 221 -82
rect 225 -86 229 -82
rect 225 -94 229 -90
rect 225 -102 229 -98
rect 225 -116 229 -106
rect 225 -124 229 -120
rect 225 -132 229 -128
rect 225 -140 229 -136
rect 233 -140 237 -82
rect 241 -86 245 -82
rect 241 -94 245 -90
rect 241 -102 245 -98
rect 241 -116 245 -106
rect 241 -124 245 -120
rect 241 -132 245 -128
rect 241 -140 245 -136
rect 249 -140 253 -82
rect 257 -86 261 -82
rect 257 -94 261 -90
rect 257 -102 261 -98
rect 257 -116 261 -106
rect 257 -124 261 -120
rect 257 -132 261 -128
rect 257 -140 261 -136
rect 265 -140 269 -82
rect 273 -86 277 -82
rect 273 -94 277 -90
rect 273 -102 277 -98
rect 273 -116 277 -106
rect 273 -124 277 -120
rect 273 -132 277 -128
rect 273 -140 277 -136
rect 281 -140 285 -82
rect 289 -86 293 -82
rect 289 -94 293 -90
rect 289 -102 293 -98
rect 289 -116 293 -106
rect 289 -124 293 -120
rect 289 -132 293 -128
rect 289 -140 293 -136
<< psubstratepcontact >>
rect 151 -184 191 -166
<< nsubstratencontact >>
rect 162 -130 191 -83
<< polysilicon >>
rect 197 -81 199 -79
rect 214 -80 288 -77
rect 214 -81 216 -80
rect 222 -81 224 -80
rect 230 -81 232 -80
rect 238 -81 240 -80
rect 246 -81 248 -80
rect 254 -81 256 -80
rect 262 -81 264 -80
rect 270 -81 272 -80
rect 278 -81 280 -80
rect 286 -81 288 -80
rect 163 -135 165 -133
rect 168 -135 170 -133
rect 177 -135 179 -133
rect 163 -149 165 -141
rect 168 -142 170 -141
rect 168 -143 174 -142
rect 168 -147 169 -143
rect 173 -147 174 -143
rect 168 -148 174 -147
rect 158 -150 165 -149
rect 158 -154 159 -150
rect 163 -154 165 -150
rect 158 -155 165 -154
rect 163 -156 165 -155
rect 171 -156 173 -148
rect 177 -149 179 -141
rect 197 -142 199 -141
rect 214 -142 216 -141
rect 222 -142 224 -141
rect 230 -142 232 -141
rect 238 -142 240 -141
rect 246 -142 248 -141
rect 254 -142 256 -141
rect 262 -142 264 -141
rect 270 -142 272 -141
rect 278 -142 280 -141
rect 286 -142 288 -141
rect 193 -147 199 -142
rect 177 -150 183 -149
rect 177 -154 178 -150
rect 182 -154 183 -150
rect 177 -155 183 -154
rect 193 -151 194 -147
rect 198 -151 199 -147
rect 193 -155 199 -151
rect 210 -143 294 -142
rect 210 -154 211 -143
rect 215 -154 294 -143
rect 210 -155 294 -154
rect 179 -156 181 -155
rect 197 -156 199 -155
rect 214 -156 216 -155
rect 222 -156 224 -155
rect 230 -156 232 -155
rect 238 -156 240 -155
rect 246 -156 248 -155
rect 254 -156 256 -155
rect 262 -156 264 -155
rect 270 -156 272 -155
rect 278 -156 280 -155
rect 286 -156 288 -155
rect 163 -164 165 -162
rect 171 -164 173 -162
rect 179 -164 181 -162
rect 197 -188 199 -186
rect 214 -187 216 -186
rect 222 -187 224 -186
rect 230 -187 232 -186
rect 238 -187 240 -186
rect 246 -187 248 -186
rect 254 -187 256 -186
rect 262 -187 264 -186
rect 270 -187 272 -186
rect 278 -187 280 -186
rect 286 -187 288 -186
rect 214 -191 288 -187
<< polycontact >>
rect 169 -147 173 -143
rect 159 -154 163 -150
rect 178 -154 182 -150
rect 194 -151 198 -147
rect 211 -154 215 -143
<< metal1 >>
rect 150 -83 192 -82
rect 150 -130 162 -83
rect 191 -130 192 -83
rect 150 -133 192 -130
rect 150 -140 155 -133
rect 171 -136 175 -133
rect 184 -140 189 -136
rect 204 -140 205 -82
rect 221 -140 222 -82
rect 237 -140 238 -82
rect 253 -140 254 -82
rect 269 -140 270 -82
rect 285 -140 286 -82
rect 150 -147 169 -143
rect 185 -147 189 -140
rect 200 -143 205 -140
rect 218 -143 222 -140
rect 234 -143 238 -140
rect 250 -143 254 -140
rect 266 -143 270 -140
rect 282 -143 286 -140
rect 200 -144 211 -143
rect 150 -154 159 -150
rect 176 -151 178 -150
rect 166 -153 178 -151
rect 170 -154 178 -153
rect 185 -151 194 -147
rect 185 -157 189 -151
rect 201 -154 211 -144
rect 218 -154 300 -143
rect 200 -157 205 -154
rect 218 -157 222 -154
rect 234 -157 238 -154
rect 250 -157 254 -154
rect 266 -157 270 -154
rect 282 -157 286 -154
rect 150 -161 158 -157
rect 166 -161 170 -157
rect 186 -161 189 -157
rect 150 -164 162 -161
rect 174 -164 178 -161
rect 150 -166 192 -164
rect 150 -184 151 -166
rect 191 -184 192 -166
rect 150 -185 192 -184
rect 204 -185 205 -157
rect 221 -185 222 -157
rect 237 -185 238 -157
rect 253 -185 254 -157
rect 269 -185 270 -157
rect 285 -185 286 -157
<< m2contact >>
rect 192 -90 196 -86
rect 192 -98 196 -94
rect 192 -106 196 -102
rect 192 -120 196 -116
rect 192 -128 196 -124
rect 192 -136 196 -132
rect 162 -140 166 -136
rect 209 -90 213 -86
rect 209 -98 213 -94
rect 209 -106 213 -102
rect 209 -120 213 -116
rect 209 -128 213 -124
rect 209 -136 213 -132
rect 225 -90 229 -86
rect 225 -98 229 -94
rect 225 -106 229 -102
rect 225 -120 229 -116
rect 225 -128 229 -124
rect 225 -136 229 -132
rect 241 -90 245 -86
rect 241 -98 245 -94
rect 241 -106 245 -102
rect 241 -120 245 -116
rect 241 -128 245 -124
rect 241 -136 245 -132
rect 257 -90 261 -86
rect 257 -98 261 -94
rect 257 -106 261 -102
rect 257 -120 261 -116
rect 257 -128 261 -124
rect 257 -136 261 -132
rect 273 -90 277 -86
rect 273 -98 277 -94
rect 273 -106 277 -102
rect 273 -120 277 -116
rect 273 -128 277 -124
rect 273 -136 277 -132
rect 289 -90 293 -86
rect 289 -98 293 -94
rect 289 -106 293 -102
rect 289 -120 293 -116
rect 289 -128 293 -124
rect 289 -136 293 -132
rect 166 -157 170 -153
rect 192 -165 196 -161
rect 192 -173 196 -169
rect 192 -181 196 -177
rect 209 -165 213 -161
rect 209 -173 213 -169
rect 209 -181 213 -177
rect 225 -165 229 -161
rect 225 -173 229 -169
rect 225 -181 229 -177
rect 241 -165 245 -161
rect 241 -173 245 -169
rect 241 -181 245 -177
rect 257 -165 261 -161
rect 257 -173 261 -169
rect 257 -181 261 -177
rect 273 -165 277 -161
rect 273 -173 277 -169
rect 273 -181 277 -177
rect 289 -165 293 -161
rect 289 -173 293 -169
rect 289 -181 293 -177
<< metal2 >>
rect 192 -86 293 -82
rect 196 -90 209 -86
rect 213 -90 225 -86
rect 229 -90 241 -86
rect 245 -90 257 -86
rect 261 -90 273 -86
rect 277 -90 289 -86
rect 192 -94 293 -90
rect 196 -98 209 -94
rect 213 -98 225 -94
rect 229 -98 241 -94
rect 245 -98 257 -94
rect 261 -98 273 -94
rect 277 -98 289 -94
rect 192 -102 293 -98
rect 196 -106 209 -102
rect 213 -106 225 -102
rect 229 -106 241 -102
rect 245 -106 257 -102
rect 261 -106 273 -102
rect 277 -106 289 -102
rect 192 -116 293 -106
rect 196 -120 209 -116
rect 213 -120 225 -116
rect 229 -120 241 -116
rect 245 -120 257 -116
rect 261 -120 273 -116
rect 277 -120 289 -116
rect 192 -124 293 -120
rect 196 -128 209 -124
rect 213 -128 225 -124
rect 229 -128 241 -124
rect 245 -128 257 -124
rect 261 -128 273 -124
rect 277 -128 289 -124
rect 192 -132 293 -128
rect 196 -136 209 -132
rect 213 -136 225 -132
rect 229 -136 241 -132
rect 245 -136 257 -132
rect 261 -136 273 -132
rect 277 -136 289 -132
rect 158 -147 162 -136
rect 192 -140 293 -136
rect 158 -151 170 -147
rect 166 -153 170 -151
rect 166 -161 170 -157
rect 192 -161 293 -157
rect 196 -165 209 -161
rect 213 -165 225 -161
rect 229 -165 241 -161
rect 245 -165 257 -161
rect 261 -165 273 -161
rect 277 -165 289 -161
rect 192 -169 293 -165
rect 196 -173 209 -169
rect 213 -173 225 -169
rect 229 -173 241 -169
rect 245 -173 257 -169
rect 261 -173 273 -169
rect 277 -173 289 -169
rect 192 -177 293 -173
rect 196 -181 209 -177
rect 213 -181 225 -177
rect 229 -181 241 -177
rect 245 -181 257 -177
rect 261 -181 273 -177
rect 277 -181 289 -177
rect 192 -185 293 -181
<< labels >>
rlabel metal1 155 -161 158 -157 1 Gnd
rlabel metal1 155 -154 159 -150 1 B
rlabel metal1 155 -147 169 -143 1 A
rlabel metal1 150 -140 155 -136 3 Vdd
rlabel metal1 218 -154 300 -143 1 Z
<< end >>
