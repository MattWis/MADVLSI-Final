magic
tech scmos
timestamp 1418787195
<< metal1 >>
rect -94 497 -57 500
rect -53 497 81 500
rect 85 497 133 500
rect 137 497 155 500
rect 111 490 155 493
rect 111 488 115 490
rect -38 474 0 478
rect 130 474 133 478
rect -94 467 -42 471
rect -87 437 -84 467
rect -31 462 0 466
rect 130 462 147 466
rect -59 450 -57 453
rect -24 450 0 454
rect 130 450 140 454
rect -87 433 -81 437
rect -59 433 -21 437
rect 111 429 155 432
rect 111 427 115 429
rect -59 417 -49 420
rect -38 413 0 417
rect 130 413 133 417
rect -31 401 0 405
rect 130 401 147 405
rect -3 389 0 393
rect 130 389 140 393
rect 111 368 155 371
rect 111 366 115 368
rect -38 352 0 356
rect 130 352 133 356
rect -94 345 -35 349
rect -87 315 -84 345
rect -10 340 0 344
rect 130 340 147 344
rect -59 328 -57 331
rect -24 328 0 332
rect 130 328 140 332
rect -87 311 -81 315
rect -59 311 -14 315
rect 111 307 155 310
rect 111 305 115 307
rect -59 295 -49 298
rect -38 291 0 295
rect 130 291 133 295
rect -10 279 0 283
rect 130 279 147 283
rect -3 267 0 271
rect 111 246 155 249
rect 111 244 115 246
rect -94 227 -28 231
rect -17 230 0 234
rect 130 230 133 234
rect -87 193 -84 227
rect -31 218 0 222
rect 130 218 147 222
rect -59 206 -57 209
rect -24 206 0 210
rect 130 206 140 210
rect -87 189 -81 193
rect -59 189 -7 193
rect 111 185 155 188
rect 111 183 115 185
rect -59 173 -49 176
rect -17 169 0 173
rect 130 169 133 173
rect -31 157 0 161
rect 130 157 147 161
rect -3 145 0 149
rect 130 145 140 149
rect 111 124 155 127
rect 111 122 115 124
rect -17 108 0 112
rect 130 108 133 112
rect -10 96 0 100
rect 130 96 147 100
rect -24 84 0 88
rect 130 84 140 88
rect 111 63 155 66
rect 111 61 115 63
rect -17 47 0 51
rect 130 47 133 51
rect -10 35 0 39
rect 130 35 147 39
rect -3 23 0 27
rect 130 23 140 27
rect -94 -7 -49 -4
rect -45 -7 88 -4
rect 92 -7 140 -4
rect 144 -7 155 -4
<< m2contact >>
rect -57 496 -53 500
rect 81 496 85 500
rect 133 496 137 500
rect -42 474 -38 478
rect 133 474 137 478
rect -42 467 -38 471
rect -35 462 -31 466
rect 147 462 151 466
rect -57 449 -53 453
rect -28 450 -24 454
rect 140 450 144 454
rect -21 433 -17 437
rect -49 416 -45 420
rect -42 413 -38 417
rect 133 413 137 417
rect -35 401 -31 405
rect 147 401 151 405
rect -7 389 -3 393
rect 140 389 144 393
rect -42 352 -38 356
rect 133 352 137 356
rect -35 345 -31 349
rect -14 340 -10 344
rect 147 340 151 344
rect -57 327 -53 331
rect -28 328 -24 332
rect 140 328 144 332
rect -14 311 -10 315
rect -49 294 -45 298
rect -42 291 -38 295
rect 133 291 137 295
rect -14 279 -10 283
rect 147 279 151 283
rect -7 267 -3 271
rect 140 267 144 271
rect -28 227 -24 231
rect -21 230 -17 234
rect 133 230 137 234
rect -35 218 -31 222
rect 147 218 151 222
rect -57 205 -53 209
rect -28 206 -24 210
rect 140 206 144 210
rect -7 189 -3 193
rect -49 172 -45 176
rect -21 169 -17 173
rect 133 169 137 173
rect -35 157 -31 161
rect 147 157 151 161
rect -7 145 -3 149
rect 140 145 144 149
rect -21 108 -17 112
rect 133 108 137 112
rect -14 96 -10 100
rect 147 96 151 100
rect -28 84 -24 88
rect 140 84 144 88
rect -21 47 -17 51
rect 133 47 137 51
rect -14 35 -10 39
rect 147 35 151 39
rect -7 23 -3 27
rect 140 23 144 27
rect -49 -7 -45 -3
rect 88 -7 92 -3
rect 140 -7 144 -3
<< metal2 >>
rect -57 453 -53 496
rect 81 488 85 496
rect -57 331 -53 449
rect -57 209 -53 327
rect -57 0 -53 205
rect -49 420 -45 488
rect -49 298 -45 416
rect -49 176 -45 294
rect -49 -3 -45 172
rect -42 478 -38 488
rect -42 471 -38 474
rect -42 417 -38 467
rect -42 356 -38 413
rect -42 295 -38 352
rect -42 0 -38 291
rect -35 466 -31 488
rect -35 405 -31 462
rect -35 349 -31 401
rect -35 222 -31 345
rect -35 161 -31 218
rect -35 0 -31 157
rect -28 454 -24 488
rect -28 332 -24 450
rect -28 231 -24 328
rect -28 210 -24 227
rect -28 88 -24 206
rect -28 0 -24 84
rect -21 437 -17 488
rect -21 234 -17 433
rect -21 173 -17 230
rect -21 112 -17 169
rect -21 51 -17 108
rect -21 0 -17 47
rect -14 344 -10 488
rect -14 315 -10 340
rect -14 283 -10 311
rect -14 100 -10 279
rect -14 39 -10 96
rect -14 0 -10 35
rect -7 393 -3 488
rect -7 271 -3 389
rect -7 193 -3 267
rect -7 149 -3 189
rect -7 27 -3 145
rect -7 0 -3 23
rect 133 478 137 496
rect 133 417 137 474
rect 133 356 137 413
rect 133 295 137 352
rect 133 234 137 291
rect 133 173 137 230
rect 133 112 137 169
rect 133 51 137 108
rect 133 0 137 47
rect 140 454 144 488
rect 140 393 144 450
rect 140 332 144 389
rect 140 271 144 328
rect 140 210 144 267
rect 140 149 144 206
rect 140 88 144 145
rect 140 27 144 84
rect 88 -3 92 0
rect 140 -3 144 23
rect 147 466 151 488
rect 147 405 151 462
rect 147 344 151 401
rect 147 283 151 340
rect 147 222 151 279
rect 147 161 151 218
rect 147 100 151 157
rect 147 39 151 96
rect 147 15 151 35
rect 147 11 155 15
rect 147 0 151 11
use inverter  inverter_0
timestamp 1418784353
transform 1 0 -80 0 1 442
box -1 -33 21 19
use 3AND  3AND_7
timestamp 1418282175
transform 1 0 65 0 1 454
box -65 -27 33 34
use PassGate  PassGate_7
timestamp 1418276510
transform 1 0 115 0 1 457
box -17 -17 15 31
use 3AND  3AND_6
timestamp 1418282175
transform 1 0 65 0 1 393
box -65 -27 33 34
use PassGate  PassGate_6
timestamp 1418276510
transform 1 0 115 0 1 396
box -17 -17 15 31
use inverter  inverter_1
timestamp 1418784353
transform 1 0 -80 0 1 320
box -1 -33 21 19
use 3AND  3AND_5
timestamp 1418282175
transform 1 0 65 0 1 332
box -65 -27 33 34
use PassGate  PassGate_5
timestamp 1418276510
transform 1 0 115 0 1 335
box -17 -17 15 31
use 3AND  3AND_4
timestamp 1418282175
transform 1 0 65 0 1 271
box -65 -27 33 34
use PassGate  PassGate_4
timestamp 1418276510
transform 1 0 115 0 1 274
box -17 -17 15 31
use inverter  inverter_2
timestamp 1418784353
transform 1 0 -80 0 1 198
box -1 -33 21 19
use 3AND  3AND_3
timestamp 1418282175
transform 1 0 65 0 1 210
box -65 -27 33 34
use PassGate  PassGate_3
timestamp 1418276510
transform 1 0 115 0 1 213
box -17 -17 15 31
use 3AND  3AND_2
timestamp 1418282175
transform 1 0 65 0 1 149
box -65 -27 33 34
use PassGate  PassGate_2
timestamp 1418276510
transform 1 0 115 0 1 152
box -17 -17 15 31
use 3AND  3AND_1
timestamp 1418282175
transform 1 0 65 0 1 88
box -65 -27 33 34
use PassGate  PassGate_1
timestamp 1418276510
transform 1 0 115 0 1 91
box -17 -17 15 31
use 3AND  3AND_0
timestamp 1418282175
transform 1 0 65 0 1 27
box -65 -27 33 34
use PassGate  PassGate_0
timestamp 1418276510
transform 1 0 115 0 1 30
box -17 -17 15 31
<< labels >>
rlabel metal2 -42 486 -38 488 4 A
rlabel metal2 -35 486 -31 488 5 B
rlabel metal2 -28 486 -24 488 5 C
rlabel metal2 -14 486 -10 488 5 Bnot
rlabel metal2 -7 486 -3 488 5 Cnot
rlabel metal2 -21 486 -17 488 5 Anot
rlabel metal1 153 63 155 66 7 bit0Input
rlabel metal1 153 124 155 127 7 bit1Input
rlabel metal1 153 185 155 188 7 bit2Input
rlabel metal1 153 246 155 249 7 bit3Input
rlabel metal1 153 307 155 310 7 bit4Input
rlabel metal1 153 368 155 371 7 bit5Input
rlabel metal1 153 429 155 432 7 bit6Input
rlabel metal1 153 490 155 493 7 bit7Input
rlabel metal1 -94 227 -92 231 1 DAC_C
rlabel metal1 -94 345 -92 349 1 DAC_B
rlabel metal1 -94 467 -92 471 1 DAC_A
rlabel metal1 -94 -7 -92 -4 1 gnd
rlabel metal1 -94 497 -92 500 4 vdd
rlabel metal1 153 497 155 500 6 Vdd
rlabel metal1 153 -7 155 -4 8 gnd
rlabel metal2 153 11 155 15 7 output
<< end >>
