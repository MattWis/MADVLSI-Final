magic
tech scmos
timestamp 1418747290
<< error_s >>
rect 796 4679 797 4683
rect 802 4679 803 4683
rect 808 4679 809 4683
rect 814 4679 815 4683
rect 820 4679 821 4683
rect 826 4679 827 4683
rect 858 4679 859 4683
rect 864 4679 865 4683
rect 870 4679 871 4683
rect 876 4679 877 4683
rect 882 4679 883 4683
rect 888 4679 889 4683
rect 1270 4679 1271 4683
rect 1276 4679 1277 4683
rect 1282 4679 1283 4683
rect 1288 4679 1289 4683
rect 1294 4679 1295 4683
rect 1300 4679 1301 4683
rect 1332 4679 1333 4683
rect 1338 4679 1339 4683
rect 1344 4679 1345 4683
rect 1350 4679 1351 4683
rect 1356 4679 1357 4683
rect 1362 4679 1363 4683
rect 1744 4679 1745 4683
rect 1750 4679 1751 4683
rect 1756 4679 1757 4683
rect 1762 4679 1763 4683
rect 1768 4679 1769 4683
rect 1774 4679 1775 4683
rect 796 4667 797 4671
rect 802 4667 803 4671
rect 808 4667 809 4671
rect 814 4667 815 4671
rect 820 4667 821 4671
rect 826 4667 827 4671
rect 858 4667 859 4671
rect 864 4667 865 4671
rect 870 4667 871 4671
rect 876 4667 877 4671
rect 882 4667 883 4671
rect 888 4667 889 4671
rect 1270 4667 1271 4671
rect 1276 4667 1277 4671
rect 1282 4667 1283 4671
rect 1288 4667 1289 4671
rect 1294 4667 1295 4671
rect 1300 4667 1301 4671
rect 1332 4667 1333 4671
rect 1338 4667 1339 4671
rect 1344 4667 1345 4671
rect 1350 4667 1351 4671
rect 1356 4667 1357 4671
rect 1362 4667 1363 4671
rect 1744 4667 1745 4671
rect 1750 4667 1751 4671
rect 1756 4667 1757 4671
rect 1762 4667 1763 4671
rect 1768 4667 1769 4671
rect 1774 4667 1775 4671
rect 796 4655 797 4659
rect 802 4655 803 4659
rect 808 4655 809 4659
rect 814 4655 815 4659
rect 820 4655 821 4659
rect 826 4655 827 4659
rect 858 4655 859 4659
rect 864 4655 865 4659
rect 870 4655 871 4659
rect 876 4655 877 4659
rect 882 4655 883 4659
rect 888 4655 889 4659
rect 1270 4655 1271 4659
rect 1276 4655 1277 4659
rect 1282 4655 1283 4659
rect 1288 4655 1289 4659
rect 1294 4655 1295 4659
rect 1300 4655 1301 4659
rect 1332 4655 1333 4659
rect 1338 4655 1339 4659
rect 1344 4655 1345 4659
rect 1350 4655 1351 4659
rect 1356 4655 1357 4659
rect 1362 4655 1363 4659
rect 1744 4655 1745 4659
rect 1750 4655 1751 4659
rect 1756 4655 1757 4659
rect 1762 4655 1763 4659
rect 1768 4655 1769 4659
rect 1774 4655 1775 4659
rect 1019 4612 1020 4616
rect 1025 4612 1026 4616
rect 1031 4612 1032 4616
rect 1037 4612 1038 4616
rect 1043 4612 1044 4616
rect 1049 4612 1050 4616
rect 1109 4612 1110 4616
rect 1115 4612 1116 4616
rect 1121 4612 1122 4616
rect 1127 4612 1128 4616
rect 1133 4612 1134 4616
rect 1139 4612 1140 4616
rect 1493 4612 1494 4616
rect 1499 4612 1500 4616
rect 1505 4612 1506 4616
rect 1511 4612 1512 4616
rect 1517 4612 1518 4616
rect 1523 4612 1524 4616
rect 1583 4612 1584 4616
rect 1589 4612 1590 4616
rect 1595 4612 1596 4616
rect 1601 4612 1602 4616
rect 1607 4612 1608 4616
rect 1613 4612 1614 4616
rect 1967 4612 1968 4616
rect 1973 4612 1974 4616
rect 1979 4612 1980 4616
rect 1985 4612 1986 4616
rect 1991 4612 1992 4616
rect 1997 4612 1998 4616
rect 2057 4612 2058 4616
rect 2063 4612 2064 4616
rect 2069 4612 2070 4616
rect 2075 4612 2076 4616
rect 2081 4612 2082 4616
rect 2087 4612 2088 4616
rect 2915 4612 2916 4616
rect 2921 4612 2922 4616
rect 2927 4612 2928 4616
rect 2933 4612 2934 4616
rect 2939 4612 2940 4616
rect 2945 4612 2946 4616
rect 3005 4612 3006 4616
rect 3011 4612 3012 4616
rect 3017 4612 3018 4616
rect 3023 4612 3024 4616
rect 3029 4612 3030 4616
rect 3035 4612 3036 4616
rect 3389 4612 3390 4616
rect 3395 4612 3396 4616
rect 3401 4612 3402 4616
rect 3407 4612 3408 4616
rect 3413 4612 3414 4616
rect 3419 4612 3420 4616
rect 3479 4612 3480 4616
rect 3485 4612 3486 4616
rect 3491 4612 3492 4616
rect 3497 4612 3498 4616
rect 3503 4612 3504 4616
rect 3509 4612 3510 4616
rect 3863 4612 3864 4616
rect 3869 4612 3870 4616
rect 3875 4612 3876 4616
rect 3881 4612 3882 4616
rect 3887 4612 3888 4616
rect 3893 4612 3894 4616
rect 3953 4612 3954 4616
rect 3959 4612 3960 4616
rect 3965 4612 3966 4616
rect 3971 4612 3972 4616
rect 3977 4612 3978 4616
rect 3983 4612 3984 4616
rect 4337 4612 4338 4616
rect 4343 4612 4344 4616
rect 4349 4612 4350 4616
rect 4355 4612 4356 4616
rect 4361 4612 4362 4616
rect 4367 4612 4368 4616
rect 4427 4612 4428 4616
rect 4433 4612 4434 4616
rect 4439 4612 4440 4616
rect 4445 4612 4446 4616
rect 4451 4612 4452 4616
rect 4457 4612 4458 4616
rect 1019 4599 1020 4603
rect 1025 4599 1026 4603
rect 1031 4599 1032 4603
rect 1037 4599 1038 4603
rect 1043 4599 1044 4603
rect 1049 4599 1050 4603
rect 1109 4599 1110 4603
rect 1115 4599 1116 4603
rect 1121 4599 1122 4603
rect 1127 4599 1128 4603
rect 1133 4599 1134 4603
rect 1139 4599 1140 4603
rect 1493 4599 1494 4603
rect 1499 4599 1500 4603
rect 1505 4599 1506 4603
rect 1511 4599 1512 4603
rect 1517 4599 1518 4603
rect 1523 4599 1524 4603
rect 1583 4599 1584 4603
rect 1589 4599 1590 4603
rect 1595 4599 1596 4603
rect 1601 4599 1602 4603
rect 1607 4599 1608 4603
rect 1613 4599 1614 4603
rect 1967 4599 1968 4603
rect 1973 4599 1974 4603
rect 1979 4599 1980 4603
rect 1985 4599 1986 4603
rect 1991 4599 1992 4603
rect 1997 4599 1998 4603
rect 2057 4599 2058 4603
rect 2063 4599 2064 4603
rect 2069 4599 2070 4603
rect 2075 4599 2076 4603
rect 2081 4599 2082 4603
rect 2087 4599 2088 4603
rect 2915 4599 2916 4603
rect 2921 4599 2922 4603
rect 2927 4599 2928 4603
rect 2933 4599 2934 4603
rect 2939 4599 2940 4603
rect 2945 4599 2946 4603
rect 3005 4599 3006 4603
rect 3011 4599 3012 4603
rect 3017 4599 3018 4603
rect 3023 4599 3024 4603
rect 3029 4599 3030 4603
rect 3035 4599 3036 4603
rect 3389 4599 3390 4603
rect 3395 4599 3396 4603
rect 3401 4599 3402 4603
rect 3407 4599 3408 4603
rect 3413 4599 3414 4603
rect 3419 4599 3420 4603
rect 3479 4599 3480 4603
rect 3485 4599 3486 4603
rect 3491 4599 3492 4603
rect 3497 4599 3498 4603
rect 3503 4599 3504 4603
rect 3509 4599 3510 4603
rect 3863 4599 3864 4603
rect 3869 4599 3870 4603
rect 3875 4599 3876 4603
rect 3881 4599 3882 4603
rect 3887 4599 3888 4603
rect 3893 4599 3894 4603
rect 3953 4599 3954 4603
rect 3959 4599 3960 4603
rect 3965 4599 3966 4603
rect 3971 4599 3972 4603
rect 3977 4599 3978 4603
rect 3983 4599 3984 4603
rect 4337 4599 4338 4603
rect 4343 4599 4344 4603
rect 4349 4599 4350 4603
rect 4355 4599 4356 4603
rect 4361 4599 4362 4603
rect 4367 4599 4368 4603
rect 4427 4599 4428 4603
rect 4433 4599 4434 4603
rect 4439 4599 4440 4603
rect 4445 4599 4446 4603
rect 4451 4599 4452 4603
rect 4457 4599 4458 4603
rect 1020 4583 1021 4586
rect 1026 4583 1027 4586
rect 1032 4583 1033 4586
rect 1038 4583 1039 4586
rect 1120 4583 1121 4586
rect 1126 4583 1127 4586
rect 1132 4583 1133 4586
rect 1138 4583 1139 4586
rect 1494 4583 1495 4586
rect 1500 4583 1501 4586
rect 1506 4583 1507 4586
rect 1512 4583 1513 4586
rect 1594 4583 1595 4586
rect 1600 4583 1601 4586
rect 1606 4583 1607 4586
rect 1612 4583 1613 4586
rect 1968 4583 1969 4586
rect 1974 4583 1975 4586
rect 1980 4583 1981 4586
rect 1986 4583 1987 4586
rect 2068 4583 2069 4586
rect 2074 4583 2075 4586
rect 2080 4583 2081 4586
rect 2086 4583 2087 4586
rect 2916 4583 2917 4586
rect 2922 4583 2923 4586
rect 2928 4583 2929 4586
rect 2934 4583 2935 4586
rect 3016 4583 3017 4586
rect 3022 4583 3023 4586
rect 3028 4583 3029 4586
rect 3034 4583 3035 4586
rect 3390 4583 3391 4586
rect 3396 4583 3397 4586
rect 3402 4583 3403 4586
rect 3408 4583 3409 4586
rect 3490 4583 3491 4586
rect 3496 4583 3497 4586
rect 3502 4583 3503 4586
rect 3508 4583 3509 4586
rect 3864 4583 3865 4586
rect 3870 4583 3871 4586
rect 3876 4583 3877 4586
rect 3882 4583 3883 4586
rect 3964 4583 3965 4586
rect 3970 4583 3971 4586
rect 3976 4583 3977 4586
rect 3982 4583 3983 4586
rect 4338 4583 4339 4586
rect 4344 4583 4345 4586
rect 4350 4583 4351 4586
rect 4356 4583 4357 4586
rect 4438 4583 4439 4586
rect 4444 4583 4445 4586
rect 4450 4583 4451 4586
rect 4456 4583 4457 4586
rect 1014 4582 1018 4583
rect 1020 4582 1024 4583
rect 1026 4582 1030 4583
rect 1032 4582 1036 4583
rect 1038 4582 1042 4583
rect 1114 4582 1118 4583
rect 1120 4582 1124 4583
rect 1126 4582 1130 4583
rect 1132 4582 1136 4583
rect 1138 4582 1142 4583
rect 1488 4582 1492 4583
rect 1494 4582 1498 4583
rect 1500 4582 1504 4583
rect 1506 4582 1510 4583
rect 1512 4582 1516 4583
rect 1588 4582 1592 4583
rect 1594 4582 1598 4583
rect 1600 4582 1604 4583
rect 1606 4582 1610 4583
rect 1612 4582 1616 4583
rect 1962 4582 1966 4583
rect 1968 4582 1972 4583
rect 1974 4582 1978 4583
rect 1980 4582 1984 4583
rect 1986 4582 1990 4583
rect 2062 4582 2066 4583
rect 2068 4582 2072 4583
rect 2074 4582 2078 4583
rect 2080 4582 2084 4583
rect 2086 4582 2090 4583
rect 2910 4582 2914 4583
rect 2916 4582 2920 4583
rect 2922 4582 2926 4583
rect 2928 4582 2932 4583
rect 2934 4582 2938 4583
rect 3010 4582 3014 4583
rect 3016 4582 3020 4583
rect 3022 4582 3026 4583
rect 3028 4582 3032 4583
rect 3034 4582 3038 4583
rect 3384 4582 3388 4583
rect 3390 4582 3394 4583
rect 3396 4582 3400 4583
rect 3402 4582 3406 4583
rect 3408 4582 3412 4583
rect 3484 4582 3488 4583
rect 3490 4582 3494 4583
rect 3496 4582 3500 4583
rect 3502 4582 3506 4583
rect 3508 4582 3512 4583
rect 3858 4582 3862 4583
rect 3864 4582 3868 4583
rect 3870 4582 3874 4583
rect 3876 4582 3880 4583
rect 3882 4582 3886 4583
rect 3958 4582 3962 4583
rect 3964 4582 3968 4583
rect 3970 4582 3974 4583
rect 3976 4582 3980 4583
rect 3982 4582 3986 4583
rect 4332 4582 4336 4583
rect 4338 4582 4342 4583
rect 4344 4582 4348 4583
rect 4350 4582 4354 4583
rect 4356 4582 4360 4583
rect 4432 4582 4436 4583
rect 4438 4582 4442 4583
rect 4444 4582 4448 4583
rect 4450 4582 4454 4583
rect 4456 4582 4460 4583
rect 1020 4576 1021 4580
rect 1026 4576 1027 4580
rect 1032 4576 1033 4580
rect 1038 4576 1039 4580
rect 1120 4576 1121 4580
rect 1126 4576 1127 4580
rect 1132 4576 1133 4580
rect 1138 4576 1139 4580
rect 1494 4576 1495 4580
rect 1500 4576 1501 4580
rect 1506 4576 1507 4580
rect 1512 4576 1513 4580
rect 1594 4576 1595 4580
rect 1600 4576 1601 4580
rect 1606 4576 1607 4580
rect 1612 4576 1613 4580
rect 1968 4576 1969 4580
rect 1974 4576 1975 4580
rect 1980 4576 1981 4580
rect 1986 4576 1987 4580
rect 2068 4576 2069 4580
rect 2074 4576 2075 4580
rect 2080 4576 2081 4580
rect 2086 4576 2087 4580
rect 2916 4576 2917 4580
rect 2922 4576 2923 4580
rect 2928 4576 2929 4580
rect 2934 4576 2935 4580
rect 3016 4576 3017 4580
rect 3022 4576 3023 4580
rect 3028 4576 3029 4580
rect 3034 4576 3035 4580
rect 3390 4576 3391 4580
rect 3396 4576 3397 4580
rect 3402 4576 3403 4580
rect 3408 4576 3409 4580
rect 3490 4576 3491 4580
rect 3496 4576 3497 4580
rect 3502 4576 3503 4580
rect 3508 4576 3509 4580
rect 3864 4576 3865 4580
rect 3870 4576 3871 4580
rect 3876 4576 3877 4580
rect 3882 4576 3883 4580
rect 3964 4576 3965 4580
rect 3970 4576 3971 4580
rect 3976 4576 3977 4580
rect 3982 4576 3983 4580
rect 4338 4576 4339 4580
rect 4344 4576 4345 4580
rect 4350 4576 4351 4580
rect 4356 4576 4357 4580
rect 4438 4576 4439 4580
rect 4444 4576 4445 4580
rect 4450 4576 4451 4580
rect 4456 4576 4457 4580
rect 1020 4570 1021 4573
rect 1026 4570 1027 4573
rect 1032 4570 1033 4573
rect 1038 4570 1039 4573
rect 1120 4570 1121 4573
rect 1126 4570 1127 4573
rect 1132 4570 1133 4573
rect 1138 4570 1139 4573
rect 1494 4570 1495 4573
rect 1500 4570 1501 4573
rect 1506 4570 1507 4573
rect 1512 4570 1513 4573
rect 1594 4570 1595 4573
rect 1600 4570 1601 4573
rect 1606 4570 1607 4573
rect 1612 4570 1613 4573
rect 1968 4570 1969 4573
rect 1974 4570 1975 4573
rect 1980 4570 1981 4573
rect 1986 4570 1987 4573
rect 2068 4570 2069 4573
rect 2074 4570 2075 4573
rect 2080 4570 2081 4573
rect 2086 4570 2087 4573
rect 2916 4570 2917 4573
rect 2922 4570 2923 4573
rect 2928 4570 2929 4573
rect 2934 4570 2935 4573
rect 3016 4570 3017 4573
rect 3022 4570 3023 4573
rect 3028 4570 3029 4573
rect 3034 4570 3035 4573
rect 3390 4570 3391 4573
rect 3396 4570 3397 4573
rect 3402 4570 3403 4573
rect 3408 4570 3409 4573
rect 3490 4570 3491 4573
rect 3496 4570 3497 4573
rect 3502 4570 3503 4573
rect 3508 4570 3509 4573
rect 3864 4570 3865 4573
rect 3870 4570 3871 4573
rect 3876 4570 3877 4573
rect 3882 4570 3883 4573
rect 3964 4570 3965 4573
rect 3970 4570 3971 4573
rect 3976 4570 3977 4573
rect 3982 4570 3983 4573
rect 4338 4570 4339 4573
rect 4344 4570 4345 4573
rect 4350 4570 4351 4573
rect 4356 4570 4357 4573
rect 4438 4570 4439 4573
rect 4444 4570 4445 4573
rect 4450 4570 4451 4573
rect 4456 4570 4457 4573
rect 1014 4569 1018 4570
rect 1020 4569 1024 4570
rect 1026 4569 1030 4570
rect 1032 4569 1036 4570
rect 1038 4569 1042 4570
rect 1114 4569 1118 4570
rect 1120 4569 1124 4570
rect 1126 4569 1130 4570
rect 1132 4569 1136 4570
rect 1138 4569 1142 4570
rect 1488 4569 1492 4570
rect 1494 4569 1498 4570
rect 1500 4569 1504 4570
rect 1506 4569 1510 4570
rect 1512 4569 1516 4570
rect 1588 4569 1592 4570
rect 1594 4569 1598 4570
rect 1600 4569 1604 4570
rect 1606 4569 1610 4570
rect 1612 4569 1616 4570
rect 1962 4569 1966 4570
rect 1968 4569 1972 4570
rect 1974 4569 1978 4570
rect 1980 4569 1984 4570
rect 1986 4569 1990 4570
rect 2062 4569 2066 4570
rect 2068 4569 2072 4570
rect 2074 4569 2078 4570
rect 2080 4569 2084 4570
rect 2086 4569 2090 4570
rect 2910 4569 2914 4570
rect 2916 4569 2920 4570
rect 2922 4569 2926 4570
rect 2928 4569 2932 4570
rect 2934 4569 2938 4570
rect 3010 4569 3014 4570
rect 3016 4569 3020 4570
rect 3022 4569 3026 4570
rect 3028 4569 3032 4570
rect 3034 4569 3038 4570
rect 3384 4569 3388 4570
rect 3390 4569 3394 4570
rect 3396 4569 3400 4570
rect 3402 4569 3406 4570
rect 3408 4569 3412 4570
rect 3484 4569 3488 4570
rect 3490 4569 3494 4570
rect 3496 4569 3500 4570
rect 3502 4569 3506 4570
rect 3508 4569 3512 4570
rect 3858 4569 3862 4570
rect 3864 4569 3868 4570
rect 3870 4569 3874 4570
rect 3876 4569 3880 4570
rect 3882 4569 3886 4570
rect 3958 4569 3962 4570
rect 3964 4569 3968 4570
rect 3970 4569 3974 4570
rect 3976 4569 3980 4570
rect 3982 4569 3986 4570
rect 4332 4569 4336 4570
rect 4338 4569 4342 4570
rect 4344 4569 4348 4570
rect 4350 4569 4354 4570
rect 4356 4569 4360 4570
rect 4432 4569 4436 4570
rect 4438 4569 4442 4570
rect 4444 4569 4448 4570
rect 4450 4569 4454 4570
rect 4456 4569 4460 4570
rect 1020 4564 1021 4567
rect 1026 4564 1027 4567
rect 1032 4564 1033 4567
rect 1038 4564 1039 4567
rect 1120 4564 1121 4567
rect 1126 4564 1127 4567
rect 1132 4564 1133 4567
rect 1138 4564 1139 4567
rect 1494 4564 1495 4567
rect 1500 4564 1501 4567
rect 1506 4564 1507 4567
rect 1512 4564 1513 4567
rect 1594 4564 1595 4567
rect 1600 4564 1601 4567
rect 1606 4564 1607 4567
rect 1612 4564 1613 4567
rect 1968 4564 1969 4567
rect 1974 4564 1975 4567
rect 1980 4564 1981 4567
rect 1986 4564 1987 4567
rect 2068 4564 2069 4567
rect 2074 4564 2075 4567
rect 2080 4564 2081 4567
rect 2086 4564 2087 4567
rect 2916 4564 2917 4567
rect 2922 4564 2923 4567
rect 2928 4564 2929 4567
rect 2934 4564 2935 4567
rect 3016 4564 3017 4567
rect 3022 4564 3023 4567
rect 3028 4564 3029 4567
rect 3034 4564 3035 4567
rect 3390 4564 3391 4567
rect 3396 4564 3397 4567
rect 3402 4564 3403 4567
rect 3408 4564 3409 4567
rect 3490 4564 3491 4567
rect 3496 4564 3497 4567
rect 3502 4564 3503 4567
rect 3508 4564 3509 4567
rect 3864 4564 3865 4567
rect 3870 4564 3871 4567
rect 3876 4564 3877 4567
rect 3882 4564 3883 4567
rect 3964 4564 3965 4567
rect 3970 4564 3971 4567
rect 3976 4564 3977 4567
rect 3982 4564 3983 4567
rect 4338 4564 4339 4567
rect 4344 4564 4345 4567
rect 4350 4564 4351 4567
rect 4356 4564 4357 4567
rect 4438 4564 4439 4567
rect 4444 4564 4445 4567
rect 4450 4564 4451 4567
rect 4456 4564 4457 4567
rect 1014 4563 1018 4564
rect 1020 4563 1024 4564
rect 1026 4563 1030 4564
rect 1032 4563 1036 4564
rect 1038 4563 1042 4564
rect 1114 4563 1118 4564
rect 1120 4563 1124 4564
rect 1126 4563 1130 4564
rect 1132 4563 1136 4564
rect 1138 4563 1142 4564
rect 1488 4563 1492 4564
rect 1494 4563 1498 4564
rect 1500 4563 1504 4564
rect 1506 4563 1510 4564
rect 1512 4563 1516 4564
rect 1588 4563 1592 4564
rect 1594 4563 1598 4564
rect 1600 4563 1604 4564
rect 1606 4563 1610 4564
rect 1612 4563 1616 4564
rect 1962 4563 1966 4564
rect 1968 4563 1972 4564
rect 1974 4563 1978 4564
rect 1980 4563 1984 4564
rect 1986 4563 1990 4564
rect 2062 4563 2066 4564
rect 2068 4563 2072 4564
rect 2074 4563 2078 4564
rect 2080 4563 2084 4564
rect 2086 4563 2090 4564
rect 2910 4563 2914 4564
rect 2916 4563 2920 4564
rect 2922 4563 2926 4564
rect 2928 4563 2932 4564
rect 2934 4563 2938 4564
rect 3010 4563 3014 4564
rect 3016 4563 3020 4564
rect 3022 4563 3026 4564
rect 3028 4563 3032 4564
rect 3034 4563 3038 4564
rect 3384 4563 3388 4564
rect 3390 4563 3394 4564
rect 3396 4563 3400 4564
rect 3402 4563 3406 4564
rect 3408 4563 3412 4564
rect 3484 4563 3488 4564
rect 3490 4563 3494 4564
rect 3496 4563 3500 4564
rect 3502 4563 3506 4564
rect 3508 4563 3512 4564
rect 3858 4563 3862 4564
rect 3864 4563 3868 4564
rect 3870 4563 3874 4564
rect 3876 4563 3880 4564
rect 3882 4563 3886 4564
rect 3958 4563 3962 4564
rect 3964 4563 3968 4564
rect 3970 4563 3974 4564
rect 3976 4563 3980 4564
rect 3982 4563 3986 4564
rect 4332 4563 4336 4564
rect 4338 4563 4342 4564
rect 4344 4563 4348 4564
rect 4350 4563 4354 4564
rect 4356 4563 4360 4564
rect 4432 4563 4436 4564
rect 4438 4563 4442 4564
rect 4444 4563 4448 4564
rect 4450 4563 4454 4564
rect 4456 4563 4460 4564
rect 1020 4558 1021 4561
rect 1026 4558 1027 4561
rect 1032 4558 1033 4561
rect 1038 4558 1039 4561
rect 1120 4558 1121 4561
rect 1126 4558 1127 4561
rect 1132 4558 1133 4561
rect 1138 4558 1139 4561
rect 1494 4558 1495 4561
rect 1500 4558 1501 4561
rect 1506 4558 1507 4561
rect 1512 4558 1513 4561
rect 1594 4558 1595 4561
rect 1600 4558 1601 4561
rect 1606 4558 1607 4561
rect 1612 4558 1613 4561
rect 1968 4558 1969 4561
rect 1974 4558 1975 4561
rect 1980 4558 1981 4561
rect 1986 4558 1987 4561
rect 2068 4558 2069 4561
rect 2074 4558 2075 4561
rect 2080 4558 2081 4561
rect 2086 4558 2087 4561
rect 2916 4558 2917 4561
rect 2922 4558 2923 4561
rect 2928 4558 2929 4561
rect 2934 4558 2935 4561
rect 3016 4558 3017 4561
rect 3022 4558 3023 4561
rect 3028 4558 3029 4561
rect 3034 4558 3035 4561
rect 3390 4558 3391 4561
rect 3396 4558 3397 4561
rect 3402 4558 3403 4561
rect 3408 4558 3409 4561
rect 3490 4558 3491 4561
rect 3496 4558 3497 4561
rect 3502 4558 3503 4561
rect 3508 4558 3509 4561
rect 3864 4558 3865 4561
rect 3870 4558 3871 4561
rect 3876 4558 3877 4561
rect 3882 4558 3883 4561
rect 3964 4558 3965 4561
rect 3970 4558 3971 4561
rect 3976 4558 3977 4561
rect 3982 4558 3983 4561
rect 4338 4558 4339 4561
rect 4344 4558 4345 4561
rect 4350 4558 4351 4561
rect 4356 4558 4357 4561
rect 4438 4558 4439 4561
rect 4444 4558 4445 4561
rect 4450 4558 4451 4561
rect 4456 4558 4457 4561
rect 1014 4557 1018 4558
rect 1020 4557 1024 4558
rect 1026 4557 1030 4558
rect 1032 4557 1036 4558
rect 1038 4557 1042 4558
rect 1114 4557 1118 4558
rect 1120 4557 1124 4558
rect 1126 4557 1130 4558
rect 1132 4557 1136 4558
rect 1138 4557 1142 4558
rect 1488 4557 1492 4558
rect 1494 4557 1498 4558
rect 1500 4557 1504 4558
rect 1506 4557 1510 4558
rect 1512 4557 1516 4558
rect 1588 4557 1592 4558
rect 1594 4557 1598 4558
rect 1600 4557 1604 4558
rect 1606 4557 1610 4558
rect 1612 4557 1616 4558
rect 1962 4557 1966 4558
rect 1968 4557 1972 4558
rect 1974 4557 1978 4558
rect 1980 4557 1984 4558
rect 1986 4557 1990 4558
rect 2062 4557 2066 4558
rect 2068 4557 2072 4558
rect 2074 4557 2078 4558
rect 2080 4557 2084 4558
rect 2086 4557 2090 4558
rect 2910 4557 2914 4558
rect 2916 4557 2920 4558
rect 2922 4557 2926 4558
rect 2928 4557 2932 4558
rect 2934 4557 2938 4558
rect 3010 4557 3014 4558
rect 3016 4557 3020 4558
rect 3022 4557 3026 4558
rect 3028 4557 3032 4558
rect 3034 4557 3038 4558
rect 3384 4557 3388 4558
rect 3390 4557 3394 4558
rect 3396 4557 3400 4558
rect 3402 4557 3406 4558
rect 3408 4557 3412 4558
rect 3484 4557 3488 4558
rect 3490 4557 3494 4558
rect 3496 4557 3500 4558
rect 3502 4557 3506 4558
rect 3508 4557 3512 4558
rect 3858 4557 3862 4558
rect 3864 4557 3868 4558
rect 3870 4557 3874 4558
rect 3876 4557 3880 4558
rect 3882 4557 3886 4558
rect 3958 4557 3962 4558
rect 3964 4557 3968 4558
rect 3970 4557 3974 4558
rect 3976 4557 3980 4558
rect 3982 4557 3986 4558
rect 4332 4557 4336 4558
rect 4338 4557 4342 4558
rect 4344 4557 4348 4558
rect 4350 4557 4354 4558
rect 4356 4557 4360 4558
rect 4432 4557 4436 4558
rect 4438 4557 4442 4558
rect 4444 4557 4448 4558
rect 4450 4557 4454 4558
rect 4456 4557 4460 4558
rect 1020 4551 1021 4555
rect 1026 4551 1027 4555
rect 1032 4551 1033 4555
rect 1038 4551 1039 4555
rect 1120 4551 1121 4555
rect 1126 4551 1127 4555
rect 1132 4551 1133 4555
rect 1138 4551 1139 4555
rect 1494 4551 1495 4555
rect 1500 4551 1501 4555
rect 1506 4551 1507 4555
rect 1512 4551 1513 4555
rect 1594 4551 1595 4555
rect 1600 4551 1601 4555
rect 1606 4551 1607 4555
rect 1612 4551 1613 4555
rect 1968 4551 1969 4555
rect 1974 4551 1975 4555
rect 1980 4551 1981 4555
rect 1986 4551 1987 4555
rect 2068 4551 2069 4555
rect 2074 4551 2075 4555
rect 2080 4551 2081 4555
rect 2086 4551 2087 4555
rect 2916 4551 2917 4555
rect 2922 4551 2923 4555
rect 2928 4551 2929 4555
rect 2934 4551 2935 4555
rect 3016 4551 3017 4555
rect 3022 4551 3023 4555
rect 3028 4551 3029 4555
rect 3034 4551 3035 4555
rect 3390 4551 3391 4555
rect 3396 4551 3397 4555
rect 3402 4551 3403 4555
rect 3408 4551 3409 4555
rect 3490 4551 3491 4555
rect 3496 4551 3497 4555
rect 3502 4551 3503 4555
rect 3508 4551 3509 4555
rect 3864 4551 3865 4555
rect 3870 4551 3871 4555
rect 3876 4551 3877 4555
rect 3882 4551 3883 4555
rect 3964 4551 3965 4555
rect 3970 4551 3971 4555
rect 3976 4551 3977 4555
rect 3982 4551 3983 4555
rect 4338 4551 4339 4555
rect 4344 4551 4345 4555
rect 4350 4551 4351 4555
rect 4356 4551 4357 4555
rect 4438 4551 4439 4555
rect 4444 4551 4445 4555
rect 4450 4551 4451 4555
rect 4456 4551 4457 4555
rect 1019 4525 1020 4529
rect 1025 4525 1026 4529
rect 1031 4525 1032 4529
rect 1037 4525 1038 4529
rect 1043 4525 1044 4529
rect 1049 4525 1050 4529
rect 1109 4525 1110 4529
rect 1115 4525 1116 4529
rect 1121 4525 1122 4529
rect 1127 4525 1128 4529
rect 1133 4525 1134 4529
rect 1139 4525 1140 4529
rect 1493 4525 1494 4529
rect 1499 4525 1500 4529
rect 1505 4525 1506 4529
rect 1511 4525 1512 4529
rect 1517 4525 1518 4529
rect 1523 4525 1524 4529
rect 1583 4525 1584 4529
rect 1589 4525 1590 4529
rect 1595 4525 1596 4529
rect 1601 4525 1602 4529
rect 1607 4525 1608 4529
rect 1613 4525 1614 4529
rect 1967 4525 1968 4529
rect 1973 4525 1974 4529
rect 1979 4525 1980 4529
rect 1985 4525 1986 4529
rect 1991 4525 1992 4529
rect 1997 4525 1998 4529
rect 2057 4525 2058 4529
rect 2063 4525 2064 4529
rect 2069 4525 2070 4529
rect 2075 4525 2076 4529
rect 2081 4525 2082 4529
rect 2087 4525 2088 4529
rect 2915 4525 2916 4529
rect 2921 4525 2922 4529
rect 2927 4525 2928 4529
rect 2933 4525 2934 4529
rect 2939 4525 2940 4529
rect 2945 4525 2946 4529
rect 3005 4525 3006 4529
rect 3011 4525 3012 4529
rect 3017 4525 3018 4529
rect 3023 4525 3024 4529
rect 3029 4525 3030 4529
rect 3035 4525 3036 4529
rect 3389 4525 3390 4529
rect 3395 4525 3396 4529
rect 3401 4525 3402 4529
rect 3407 4525 3408 4529
rect 3413 4525 3414 4529
rect 3419 4525 3420 4529
rect 3479 4525 3480 4529
rect 3485 4525 3486 4529
rect 3491 4525 3492 4529
rect 3497 4525 3498 4529
rect 3503 4525 3504 4529
rect 3509 4525 3510 4529
rect 3863 4525 3864 4529
rect 3869 4525 3870 4529
rect 3875 4525 3876 4529
rect 3881 4525 3882 4529
rect 3887 4525 3888 4529
rect 3893 4525 3894 4529
rect 3953 4525 3954 4529
rect 3959 4525 3960 4529
rect 3965 4525 3966 4529
rect 3971 4525 3972 4529
rect 3977 4525 3978 4529
rect 3983 4525 3984 4529
rect 4337 4525 4338 4529
rect 4343 4525 4344 4529
rect 4349 4525 4350 4529
rect 4355 4525 4356 4529
rect 4361 4525 4362 4529
rect 4367 4525 4368 4529
rect 4427 4525 4428 4529
rect 4433 4525 4434 4529
rect 4439 4525 4440 4529
rect 4445 4525 4446 4529
rect 4451 4525 4452 4529
rect 4457 4525 4458 4529
rect 1019 4507 1020 4511
rect 1025 4507 1026 4511
rect 1031 4507 1032 4511
rect 1037 4507 1038 4511
rect 1043 4507 1044 4511
rect 1049 4507 1050 4511
rect 1109 4507 1110 4511
rect 1115 4507 1116 4511
rect 1121 4507 1122 4511
rect 1127 4507 1128 4511
rect 1133 4507 1134 4511
rect 1139 4507 1140 4511
rect 1493 4507 1494 4511
rect 1499 4507 1500 4511
rect 1505 4507 1506 4511
rect 1511 4507 1512 4511
rect 1517 4507 1518 4511
rect 1523 4507 1524 4511
rect 1583 4507 1584 4511
rect 1589 4507 1590 4511
rect 1595 4507 1596 4511
rect 1601 4507 1602 4511
rect 1607 4507 1608 4511
rect 1613 4507 1614 4511
rect 1967 4507 1968 4511
rect 1973 4507 1974 4511
rect 1979 4507 1980 4511
rect 1985 4507 1986 4511
rect 1991 4507 1992 4511
rect 1997 4507 1998 4511
rect 2057 4507 2058 4511
rect 2063 4507 2064 4511
rect 2069 4507 2070 4511
rect 2075 4507 2076 4511
rect 2081 4507 2082 4511
rect 2087 4507 2088 4511
rect 2915 4507 2916 4511
rect 2921 4507 2922 4511
rect 2927 4507 2928 4511
rect 2933 4507 2934 4511
rect 2939 4507 2940 4511
rect 2945 4507 2946 4511
rect 3005 4507 3006 4511
rect 3011 4507 3012 4511
rect 3017 4507 3018 4511
rect 3023 4507 3024 4511
rect 3029 4507 3030 4511
rect 3035 4507 3036 4511
rect 3389 4507 3390 4511
rect 3395 4507 3396 4511
rect 3401 4507 3402 4511
rect 3407 4507 3408 4511
rect 3413 4507 3414 4511
rect 3419 4507 3420 4511
rect 3479 4507 3480 4511
rect 3485 4507 3486 4511
rect 3491 4507 3492 4511
rect 3497 4507 3498 4511
rect 3503 4507 3504 4511
rect 3509 4507 3510 4511
rect 3863 4507 3864 4511
rect 3869 4507 3870 4511
rect 3875 4507 3876 4511
rect 3881 4507 3882 4511
rect 3887 4507 3888 4511
rect 3893 4507 3894 4511
rect 3953 4507 3954 4511
rect 3959 4507 3960 4511
rect 3965 4507 3966 4511
rect 3971 4507 3972 4511
rect 3977 4507 3978 4511
rect 3983 4507 3984 4511
rect 4337 4507 4338 4511
rect 4343 4507 4344 4511
rect 4349 4507 4350 4511
rect 4355 4507 4356 4511
rect 4361 4507 4362 4511
rect 4367 4507 4368 4511
rect 4427 4507 4428 4511
rect 4433 4507 4434 4511
rect 4439 4507 4440 4511
rect 4445 4507 4446 4511
rect 4451 4507 4452 4511
rect 4457 4507 4458 4511
rect 4507 4457 4511 4458
rect 4525 4457 4529 4458
rect 4557 4457 4558 4460
rect 4563 4457 4564 4460
rect 4569 4457 4570 4460
rect 4582 4457 4583 4460
rect 4599 4457 4603 4458
rect 4612 4457 4616 4458
rect 4551 4456 4555 4457
rect 4557 4456 4561 4457
rect 4563 4456 4567 4457
rect 4569 4456 4573 4457
rect 4576 4456 4580 4457
rect 4582 4456 4586 4457
rect 4507 4451 4511 4452
rect 4525 4451 4529 4452
rect 4557 4451 4558 4454
rect 4563 4451 4564 4454
rect 4569 4451 4570 4454
rect 4582 4451 4583 4454
rect 4599 4451 4603 4452
rect 4612 4451 4616 4452
rect 4551 4450 4555 4451
rect 4557 4450 4561 4451
rect 4563 4450 4567 4451
rect 4569 4450 4573 4451
rect 4576 4450 4580 4451
rect 4582 4450 4586 4451
rect 4507 4445 4511 4446
rect 4525 4445 4529 4446
rect 4557 4445 4558 4448
rect 4563 4445 4564 4448
rect 4569 4445 4570 4448
rect 4582 4445 4583 4448
rect 4599 4445 4603 4446
rect 4612 4445 4616 4446
rect 4551 4444 4555 4445
rect 4557 4444 4561 4445
rect 4563 4444 4567 4445
rect 4569 4444 4573 4445
rect 4576 4444 4580 4445
rect 4582 4444 4586 4445
rect 4507 4439 4511 4440
rect 4525 4439 4529 4440
rect 4557 4439 4558 4442
rect 4563 4439 4564 4442
rect 4569 4439 4570 4442
rect 4582 4439 4583 4442
rect 4599 4439 4603 4440
rect 4612 4439 4616 4440
rect 4551 4438 4555 4439
rect 4557 4438 4561 4439
rect 4563 4438 4567 4439
rect 4569 4438 4573 4439
rect 4576 4438 4580 4439
rect 4582 4438 4586 4439
rect 4507 4433 4511 4434
rect 4525 4433 4529 4434
rect 4557 4432 4558 4436
rect 4563 4432 4564 4436
rect 4569 4432 4570 4436
rect 4582 4432 4583 4436
rect 4599 4433 4603 4434
rect 4612 4433 4616 4434
rect 4507 4427 4511 4428
rect 4525 4427 4529 4428
rect 4599 4427 4603 4428
rect 4612 4427 4616 4428
rect 4507 4367 4511 4368
rect 4525 4367 4529 4368
rect 4599 4367 4603 4368
rect 4612 4367 4616 4368
rect 4507 4361 4511 4362
rect 4525 4361 4529 4362
rect 4599 4361 4603 4362
rect 4612 4361 4616 4362
rect 4557 4357 4558 4360
rect 4563 4357 4564 4360
rect 4569 4357 4570 4360
rect 4582 4357 4583 4360
rect 4551 4356 4555 4357
rect 4557 4356 4561 4357
rect 4563 4356 4567 4357
rect 4569 4356 4573 4357
rect 4576 4356 4580 4357
rect 4582 4356 4586 4357
rect 4507 4355 4511 4356
rect 4525 4355 4529 4356
rect 4599 4355 4603 4356
rect 4612 4355 4616 4356
rect 4557 4351 4558 4354
rect 4563 4351 4564 4354
rect 4569 4351 4570 4354
rect 4582 4351 4583 4354
rect 4551 4350 4555 4351
rect 4557 4350 4561 4351
rect 4563 4350 4567 4351
rect 4569 4350 4573 4351
rect 4576 4350 4580 4351
rect 4582 4350 4586 4351
rect 4507 4349 4511 4350
rect 4525 4349 4529 4350
rect 4599 4349 4603 4350
rect 4612 4349 4616 4350
rect 4557 4345 4558 4348
rect 4563 4345 4564 4348
rect 4569 4345 4570 4348
rect 4582 4345 4583 4348
rect 4551 4344 4555 4345
rect 4557 4344 4561 4345
rect 4563 4344 4567 4345
rect 4569 4344 4573 4345
rect 4576 4344 4580 4345
rect 4582 4344 4586 4345
rect 4507 4343 4511 4344
rect 4525 4343 4529 4344
rect 4599 4343 4603 4344
rect 4612 4343 4616 4344
rect 4557 4339 4558 4342
rect 4563 4339 4564 4342
rect 4569 4339 4570 4342
rect 4582 4339 4583 4342
rect 4551 4338 4555 4339
rect 4557 4338 4561 4339
rect 4563 4338 4567 4339
rect 4569 4338 4573 4339
rect 4576 4338 4580 4339
rect 4582 4338 4586 4339
rect 4507 4337 4511 4338
rect 4525 4337 4529 4338
rect 4599 4337 4603 4338
rect 4612 4337 4616 4338
rect 4557 4332 4558 4336
rect 4563 4332 4564 4336
rect 4569 4332 4570 4336
rect 4582 4332 4583 4336
rect 4507 3983 4511 3984
rect 4525 3983 4529 3984
rect 4557 3983 4558 3986
rect 4563 3983 4564 3986
rect 4569 3983 4570 3986
rect 4582 3983 4583 3986
rect 4599 3983 4603 3984
rect 4612 3983 4616 3984
rect 4551 3982 4555 3983
rect 4557 3982 4561 3983
rect 4563 3982 4567 3983
rect 4569 3982 4573 3983
rect 4576 3982 4580 3983
rect 4582 3982 4586 3983
rect 4507 3977 4511 3978
rect 4525 3977 4529 3978
rect 4557 3977 4558 3980
rect 4563 3977 4564 3980
rect 4569 3977 4570 3980
rect 4582 3977 4583 3980
rect 4599 3977 4603 3978
rect 4612 3977 4616 3978
rect 4551 3976 4555 3977
rect 4557 3976 4561 3977
rect 4563 3976 4567 3977
rect 4569 3976 4573 3977
rect 4576 3976 4580 3977
rect 4582 3976 4586 3977
rect 4507 3971 4511 3972
rect 4525 3971 4529 3972
rect 4557 3971 4558 3974
rect 4563 3971 4564 3974
rect 4569 3971 4570 3974
rect 4582 3971 4583 3974
rect 4599 3971 4603 3972
rect 4612 3971 4616 3972
rect 4551 3970 4555 3971
rect 4557 3970 4561 3971
rect 4563 3970 4567 3971
rect 4569 3970 4573 3971
rect 4576 3970 4580 3971
rect 4582 3970 4586 3971
rect 4507 3965 4511 3966
rect 4525 3965 4529 3966
rect 4557 3965 4558 3968
rect 4563 3965 4564 3968
rect 4569 3965 4570 3968
rect 4582 3965 4583 3968
rect 4599 3965 4603 3966
rect 4612 3965 4616 3966
rect 4551 3964 4555 3965
rect 4557 3964 4561 3965
rect 4563 3964 4567 3965
rect 4569 3964 4573 3965
rect 4576 3964 4580 3965
rect 4582 3964 4586 3965
rect 4507 3959 4511 3960
rect 4525 3959 4529 3960
rect 4557 3958 4558 3962
rect 4563 3958 4564 3962
rect 4569 3958 4570 3962
rect 4582 3958 4583 3962
rect 4599 3959 4603 3960
rect 4612 3959 4616 3960
rect 4507 3953 4511 3954
rect 4525 3953 4529 3954
rect 4599 3953 4603 3954
rect 4612 3953 4616 3954
rect 4507 3893 4511 3894
rect 4525 3893 4529 3894
rect 4599 3893 4603 3894
rect 4612 3893 4616 3894
rect 4507 3887 4511 3888
rect 4525 3887 4529 3888
rect 4599 3887 4603 3888
rect 4612 3887 4616 3888
rect 4557 3883 4558 3886
rect 4563 3883 4564 3886
rect 4569 3883 4570 3886
rect 4582 3883 4583 3886
rect 4551 3882 4555 3883
rect 4557 3882 4561 3883
rect 4563 3882 4567 3883
rect 4569 3882 4573 3883
rect 4576 3882 4580 3883
rect 4582 3882 4586 3883
rect 4507 3881 4511 3882
rect 4525 3881 4529 3882
rect 4599 3881 4603 3882
rect 4612 3881 4616 3882
rect 4557 3877 4558 3880
rect 4563 3877 4564 3880
rect 4569 3877 4570 3880
rect 4582 3877 4583 3880
rect 4551 3876 4555 3877
rect 4557 3876 4561 3877
rect 4563 3876 4567 3877
rect 4569 3876 4573 3877
rect 4576 3876 4580 3877
rect 4582 3876 4586 3877
rect 4507 3875 4511 3876
rect 4525 3875 4529 3876
rect 4599 3875 4603 3876
rect 4612 3875 4616 3876
rect 4557 3871 4558 3874
rect 4563 3871 4564 3874
rect 4569 3871 4570 3874
rect 4582 3871 4583 3874
rect 4551 3870 4555 3871
rect 4557 3870 4561 3871
rect 4563 3870 4567 3871
rect 4569 3870 4573 3871
rect 4576 3870 4580 3871
rect 4582 3870 4586 3871
rect 4507 3869 4511 3870
rect 4525 3869 4529 3870
rect 4599 3869 4603 3870
rect 4612 3869 4616 3870
rect 4557 3865 4558 3868
rect 4563 3865 4564 3868
rect 4569 3865 4570 3868
rect 4582 3865 4583 3868
rect 4551 3864 4555 3865
rect 4557 3864 4561 3865
rect 4563 3864 4567 3865
rect 4569 3864 4573 3865
rect 4576 3864 4580 3865
rect 4582 3864 4586 3865
rect 4507 3863 4511 3864
rect 4525 3863 4529 3864
rect 4599 3863 4603 3864
rect 4612 3863 4616 3864
rect 4557 3858 4558 3862
rect 4563 3858 4564 3862
rect 4569 3858 4570 3862
rect 4582 3858 4583 3862
<< nwell >>
rect 3370 4228 3515 4378
<< polysilicon >>
rect 3215 4369 3221 4374
rect 3398 4372 3446 4373
rect 3398 4367 3399 4372
rect 3445 4367 3446 4372
rect 3398 4366 3446 4367
rect 3398 4365 3404 4366
rect 3419 4365 3425 4366
rect 3440 4365 3446 4366
rect 3808 4358 3814 4363
rect 3398 4244 3404 4245
rect 3419 4244 3425 4245
rect 3440 4244 3446 4245
rect 3398 4243 3446 4244
rect 3398 4238 3399 4243
rect 3430 4238 3446 4243
rect 3398 4237 3446 4238
<< pdiffusion >>
rect 3392 4364 3398 4365
rect 3392 4290 3393 4364
rect 3397 4290 3398 4364
rect 3392 4268 3398 4290
rect 3392 4246 3393 4268
rect 3397 4246 3398 4268
rect 3392 4245 3398 4246
rect 3404 4364 3410 4365
rect 3404 4358 3405 4364
rect 3409 4358 3410 4364
rect 3404 4354 3410 4358
rect 3404 4350 3405 4354
rect 3409 4350 3410 4354
rect 3404 4346 3410 4350
rect 3404 4342 3405 4346
rect 3409 4342 3410 4346
rect 3404 4338 3410 4342
rect 3404 4334 3405 4338
rect 3409 4334 3410 4338
rect 3404 4330 3410 4334
rect 3404 4326 3405 4330
rect 3409 4326 3410 4330
rect 3404 4322 3410 4326
rect 3404 4318 3405 4322
rect 3409 4318 3410 4322
rect 3404 4314 3410 4318
rect 3404 4310 3405 4314
rect 3409 4310 3410 4314
rect 3404 4306 3410 4310
rect 3404 4302 3405 4306
rect 3409 4302 3410 4306
rect 3404 4298 3410 4302
rect 3404 4294 3405 4298
rect 3409 4294 3410 4298
rect 3404 4290 3410 4294
rect 3404 4286 3405 4290
rect 3409 4286 3410 4290
rect 3404 4282 3410 4286
rect 3404 4278 3405 4282
rect 3409 4278 3410 4282
rect 3404 4274 3410 4278
rect 3404 4270 3405 4274
rect 3409 4270 3410 4274
rect 3404 4266 3410 4270
rect 3404 4262 3405 4266
rect 3409 4262 3410 4266
rect 3404 4258 3410 4262
rect 3404 4254 3405 4258
rect 3409 4254 3410 4258
rect 3404 4250 3410 4254
rect 3404 4246 3405 4250
rect 3409 4246 3410 4250
rect 3404 4245 3410 4246
rect 3413 4364 3419 4365
rect 3413 4246 3414 4364
rect 3418 4246 3419 4364
rect 3413 4245 3419 4246
rect 3425 4364 3431 4365
rect 3425 4358 3426 4364
rect 3430 4358 3431 4364
rect 3425 4354 3431 4358
rect 3425 4350 3426 4354
rect 3430 4350 3431 4354
rect 3425 4346 3431 4350
rect 3425 4342 3426 4346
rect 3430 4342 3431 4346
rect 3425 4338 3431 4342
rect 3425 4334 3426 4338
rect 3430 4334 3431 4338
rect 3425 4330 3431 4334
rect 3425 4326 3426 4330
rect 3430 4326 3431 4330
rect 3425 4322 3431 4326
rect 3425 4318 3426 4322
rect 3430 4318 3431 4322
rect 3425 4314 3431 4318
rect 3425 4310 3426 4314
rect 3430 4310 3431 4314
rect 3425 4306 3431 4310
rect 3425 4302 3426 4306
rect 3430 4302 3431 4306
rect 3425 4298 3431 4302
rect 3425 4294 3426 4298
rect 3430 4294 3431 4298
rect 3425 4290 3431 4294
rect 3425 4286 3426 4290
rect 3430 4286 3431 4290
rect 3425 4282 3431 4286
rect 3425 4278 3426 4282
rect 3430 4278 3431 4282
rect 3425 4274 3431 4278
rect 3425 4270 3426 4274
rect 3430 4270 3431 4274
rect 3425 4266 3431 4270
rect 3425 4262 3426 4266
rect 3430 4262 3431 4266
rect 3425 4258 3431 4262
rect 3425 4254 3426 4258
rect 3430 4254 3431 4258
rect 3425 4250 3431 4254
rect 3425 4246 3426 4250
rect 3430 4246 3431 4250
rect 3425 4245 3431 4246
rect 3434 4364 3440 4365
rect 3434 4246 3435 4364
rect 3439 4246 3440 4364
rect 3434 4245 3440 4246
rect 3446 4364 3452 4365
rect 3446 4358 3447 4364
rect 3451 4358 3452 4364
rect 3446 4354 3452 4358
rect 3446 4350 3447 4354
rect 3451 4350 3452 4354
rect 3446 4346 3452 4350
rect 3446 4342 3447 4346
rect 3451 4342 3452 4346
rect 3446 4338 3452 4342
rect 3446 4334 3447 4338
rect 3451 4334 3452 4338
rect 3446 4330 3452 4334
rect 3446 4326 3447 4330
rect 3451 4326 3452 4330
rect 3446 4322 3452 4326
rect 3446 4318 3447 4322
rect 3451 4318 3452 4322
rect 3446 4314 3452 4318
rect 3446 4310 3447 4314
rect 3451 4310 3452 4314
rect 3446 4306 3452 4310
rect 3446 4302 3447 4306
rect 3451 4302 3452 4306
rect 3446 4298 3452 4302
rect 3446 4294 3447 4298
rect 3451 4294 3452 4298
rect 3446 4290 3452 4294
rect 3446 4286 3447 4290
rect 3451 4286 3452 4290
rect 3446 4282 3452 4286
rect 3446 4278 3447 4282
rect 3451 4278 3452 4282
rect 3446 4274 3452 4278
rect 3446 4270 3447 4274
rect 3451 4270 3452 4274
rect 3446 4266 3452 4270
rect 3446 4262 3447 4266
rect 3451 4262 3452 4266
rect 3446 4258 3452 4262
rect 3446 4254 3447 4258
rect 3451 4254 3452 4258
rect 3446 4250 3452 4254
rect 3446 4246 3447 4250
rect 3451 4246 3452 4250
rect 3446 4245 3452 4246
<< metal1 >>
rect 1182 4528 1244 4529
rect 1013 4390 1053 4496
rect 1070 4404 1086 4496
rect 1159 4487 1244 4528
rect 1175 4486 1244 4487
rect 1198 4452 1244 4486
rect 1544 4474 1560 4507
rect 2018 4482 2034 4504
rect 1250 4404 1560 4474
rect 2006 4473 2047 4482
rect 1070 4393 1096 4404
rect 1244 4400 1560 4404
rect 1244 4393 1731 4397
rect 1013 4272 1101 4390
rect 1252 4381 1731 4393
rect 1289 4375 1731 4381
rect 1289 4316 1737 4375
rect 1576 3948 1737 4316
rect 1981 4056 2072 4473
rect 2865 4067 2904 4500
rect 2910 4383 2948 4502
rect 3182 4463 3200 4464
rect 3182 4462 3346 4463
rect 3440 4462 3456 4511
rect 3182 4447 3456 4462
rect 3857 4460 3897 4489
rect 2910 4357 3176 4383
rect 3182 4364 3200 4447
rect 3344 4446 3456 4447
rect 3817 4382 3897 4460
rect 3414 4364 3418 4367
rect 2910 4343 3121 4357
rect 2910 4330 3058 4343
rect 3451 4358 3507 4359
rect 3451 4250 3463 4358
rect 3817 4346 3853 4382
rect 2865 4064 3051 4067
rect 1979 4007 2838 4056
rect 2865 4034 3214 4064
rect 3236 4007 3289 4246
rect 3414 4243 3418 4246
rect 3435 4242 3439 4246
rect 3435 4234 3458 4242
rect 3914 4238 3930 4505
rect 3431 4097 3458 4234
rect 3826 4202 3930 4238
rect 3431 4095 3635 4097
rect 3431 4061 3638 4095
rect 3991 4090 4031 4494
rect 4394 4388 4492 4404
rect 4394 4164 4467 4388
rect 4199 4108 4467 4164
rect 4199 4104 4465 4108
rect 3431 4060 3635 4061
rect 3771 4051 4031 4090
rect 4200 4103 4465 4104
rect 1979 3962 3289 4007
rect 2769 3961 3289 3962
rect 1576 3947 3599 3948
rect 4200 3947 4325 4103
rect 1576 3847 4325 3947
<< metal2 >>
rect 3485 4491 3513 4492
rect 2966 4417 2982 4491
rect 2966 4400 3228 4417
rect 2966 4399 3037 4400
rect 3212 4372 3227 4400
rect 3212 4368 3216 4372
rect 3220 4368 3227 4372
rect 3212 4364 3227 4368
rect 3473 4364 3513 4491
rect 4388 4477 4404 4487
rect 3805 4387 4404 4477
rect 3405 4358 3513 4364
rect 3409 4354 3426 4358
rect 3430 4354 3447 4358
rect 3451 4354 3513 4358
rect 3806 4366 4404 4387
rect 3806 4362 3816 4366
rect 3806 4358 3809 4362
rect 3813 4358 3816 4362
rect 3806 4354 3816 4358
rect 3405 4350 3513 4354
rect 3409 4346 3426 4350
rect 3430 4346 3447 4350
rect 3451 4346 3513 4350
rect 3405 4342 3513 4346
rect 3409 4338 3426 4342
rect 3430 4338 3447 4342
rect 3451 4338 3513 4342
rect 3405 4334 3513 4338
rect 3409 4330 3426 4334
rect 3430 4330 3447 4334
rect 3451 4330 3513 4334
rect 3405 4326 3513 4330
rect 3409 4322 3426 4326
rect 3430 4322 3447 4326
rect 3451 4322 3513 4326
rect 3405 4318 3513 4322
rect 3409 4314 3426 4318
rect 3430 4314 3447 4318
rect 3451 4314 3513 4318
rect 3405 4310 3513 4314
rect 3409 4306 3426 4310
rect 3430 4306 3447 4310
rect 3451 4306 3513 4310
rect 3405 4302 3513 4306
rect 3409 4298 3426 4302
rect 3430 4298 3447 4302
rect 3451 4298 3513 4302
rect 3405 4294 3513 4298
rect 3106 4290 3395 4291
rect 3409 4290 3426 4294
rect 3430 4290 3447 4294
rect 3451 4290 3513 4294
rect 3106 4268 3393 4290
rect 3405 4286 3513 4290
rect 3409 4282 3426 4286
rect 3430 4282 3447 4286
rect 3451 4282 3513 4286
rect 3405 4278 3513 4282
rect 3409 4274 3426 4278
rect 3430 4274 3447 4278
rect 3451 4274 3513 4278
rect 3405 4270 3513 4274
rect 3106 4267 3395 4268
rect 3106 4266 3149 4267
rect 3409 4266 3426 4270
rect 3430 4266 3447 4270
rect 3451 4266 3513 4270
rect 3106 4172 3126 4266
rect 3405 4262 3513 4266
rect 3409 4258 3426 4262
rect 3430 4258 3447 4262
rect 3451 4258 3513 4262
rect 3405 4254 3513 4258
rect 3409 4250 3426 4254
rect 3430 4250 3447 4254
rect 3451 4250 3513 4254
rect 3405 4246 3513 4250
rect 3039 4159 3126 4172
rect 3039 4099 3056 4159
rect 3039 4095 3040 4099
rect 3044 4095 3056 4099
rect 3039 4092 3056 4095
<< ptransistor >>
rect 3398 4245 3404 4365
rect 3419 4245 3425 4365
rect 3440 4245 3446 4365
<< polycontact >>
rect 3399 4367 3445 4372
rect 3399 4238 3430 4243
<< pdcontact >>
rect 3393 4290 3397 4364
rect 3393 4246 3397 4268
rect 3405 4358 3409 4364
rect 3405 4350 3409 4354
rect 3405 4342 3409 4346
rect 3405 4334 3409 4338
rect 3405 4326 3409 4330
rect 3405 4318 3409 4322
rect 3405 4310 3409 4314
rect 3405 4302 3409 4306
rect 3405 4294 3409 4298
rect 3405 4286 3409 4290
rect 3405 4278 3409 4282
rect 3405 4270 3409 4274
rect 3405 4262 3409 4266
rect 3405 4254 3409 4258
rect 3405 4246 3409 4250
rect 3414 4246 3418 4364
rect 3426 4358 3430 4364
rect 3426 4350 3430 4354
rect 3426 4342 3430 4346
rect 3426 4334 3430 4338
rect 3426 4326 3430 4330
rect 3426 4318 3430 4322
rect 3426 4310 3430 4314
rect 3426 4302 3430 4306
rect 3426 4294 3430 4298
rect 3426 4286 3430 4290
rect 3426 4278 3430 4282
rect 3426 4270 3430 4274
rect 3426 4262 3430 4266
rect 3426 4254 3430 4258
rect 3426 4246 3430 4250
rect 3435 4246 3439 4364
rect 3447 4358 3451 4364
rect 3447 4350 3451 4354
rect 3447 4342 3451 4346
rect 3447 4334 3451 4338
rect 3447 4326 3451 4330
rect 3447 4318 3451 4322
rect 3447 4310 3451 4314
rect 3447 4302 3451 4306
rect 3447 4294 3451 4298
rect 3447 4286 3451 4290
rect 3447 4278 3451 4282
rect 3447 4270 3451 4274
rect 3447 4262 3451 4266
rect 3447 4254 3451 4258
rect 3447 4246 3451 4250
<< m2contact >>
rect 3216 4368 3220 4372
rect 3393 4268 3397 4290
rect 3405 4354 3409 4358
rect 3405 4346 3409 4350
rect 3405 4338 3409 4342
rect 3405 4330 3409 4334
rect 3405 4322 3409 4326
rect 3405 4314 3409 4318
rect 3405 4306 3409 4310
rect 3405 4298 3409 4302
rect 3405 4290 3409 4294
rect 3405 4282 3409 4286
rect 3405 4274 3409 4278
rect 3405 4266 3409 4270
rect 3405 4258 3409 4262
rect 3405 4250 3409 4254
rect 3426 4354 3430 4358
rect 3426 4346 3430 4350
rect 3426 4338 3430 4342
rect 3426 4330 3430 4334
rect 3426 4322 3430 4326
rect 3426 4314 3430 4318
rect 3426 4306 3430 4310
rect 3426 4298 3430 4302
rect 3426 4290 3430 4294
rect 3426 4282 3430 4286
rect 3426 4274 3430 4278
rect 3426 4266 3430 4270
rect 3426 4258 3430 4262
rect 3426 4250 3430 4254
rect 3809 4358 3813 4362
rect 3447 4354 3451 4358
rect 3447 4346 3451 4350
rect 3447 4338 3451 4342
rect 3447 4330 3451 4334
rect 3447 4322 3451 4326
rect 3447 4314 3451 4318
rect 3447 4306 3451 4310
rect 3447 4298 3451 4302
rect 3447 4290 3451 4294
rect 3447 4282 3451 4286
rect 3447 4274 3451 4278
rect 3447 4266 3451 4270
rect 3447 4258 3451 4262
rect 3447 4250 3451 4254
rect 3040 4095 3044 4099
<< nsubstratencontact >>
rect 3463 4250 3508 4358
use blankpad  blankpad_11
timestamp 1259953556
transform -1 0 841 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_0
timestamp 1259953556
transform -1 0 1315 0 -1 5000
box -2 0 476 513
use inorpad  inorpad_1
timestamp 1259953556
transform -1 0 1789 0 -1 5000
box -2 0 476 513
use inpad  inpad_9
timestamp 1259953556
transform -1 0 2263 0 -1 5000
box -2 0 476 513
use inpad  inpad_8
timestamp 1259953556
transform -1 0 2737 0 -1 5000
box -2 0 476 513
use inpad  inpad_7
timestamp 1259953556
transform -1 0 3211 0 -1 5000
box -2 0 476 513
use inpad  inpad_6
timestamp 1259953556
transform -1 0 3685 0 -1 5000
box -2 0 476 513
use inpad  inpad_5
timestamp 1259953556
transform -1 0 4159 0 -1 5000
box -2 0 476 513
use inpadp2  inpadp2_0
timestamp 1418747170
transform -1 0 4633 0 -1 5000
box -2 0 476 513
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 4487
box 0 0 5000 513
use 2-OR  2-OR_0
timestamp 1418434502
transform -1 0 1392 0 -1 4250
box 147 -223 302 -14
use blankpad  blankpad_27
timestamp 1259953556
transform 0 1 0 -1 0 4633
box -2 0 476 513
use Opamp  Opamp_0
timestamp 1418333453
transform 1 0 3221 0 1 4072
box -193 -11 77 303
use Opamp  Opamp_1
timestamp 1418333453
transform 1 0 3814 0 1 4062
box -193 -11 77 303
use inpad  inpad_3
timestamp 1259953556
transform 0 -1 5000 1 0 4159
box -2 0 476 513
use inpad  inpad_12
timestamp 1259953556
transform 0 1 0 -1 0 4159
box -2 0 476 513
use inpad  inpad_13
timestamp 1259953556
transform 0 1 0 -1 0 3685
box -2 0 476 513
use inpad  inpad_14
timestamp 1259953556
transform 0 1 0 -1 0 3211
box -2 0 476 513
use inpad  inpad_15
timestamp 1259953556
transform 0 1 0 -1 0 2737
box -2 0 476 513
use inpad  inpad_16
timestamp 1259953556
transform 0 1 0 -1 0 2263
box -2 0 476 513
use inpad  inpad_17
timestamp 1259953556
transform 0 1 0 -1 0 1789
box -2 0 476 513
use inpad  inpad_18
timestamp 1259953556
transform 0 1 0 -1 0 1315
box -2 0 476 513
use inpad  inpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 3685
box -2 0 476 513
use inpad  inpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 3211
box -2 0 476 513
use inpad  inpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 2737
box -2 0 476 513
use blankpad  blankpad_6
timestamp 1259953556
transform 0 -1 5000 1 0 2263
box -2 0 476 513
use blankpad  blankpad_7
timestamp 1259953556
transform 0 -1 5000 1 0 1789
box -2 0 476 513
use blankpad  blankpad_8
timestamp 1259953556
transform 0 -1 5000 1 0 1315
box -2 0 476 513
use blankpad  blankpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 841
box -2 0 476 513
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 367
box 2 2 513 4264
use blankpad  blankpad_29
timestamp 1259953556
transform 0 1 0 -1 0 841
box -2 0 476 513
use blankpad  blankpad_18
timestamp 1259953556
transform 1 0 367 0 1 0
box -2 0 476 513
use blankpad  blankpad_19
timestamp 1259953556
transform 1 0 841 0 1 0
box -2 0 476 513
use blankpad  blankpad_26
timestamp 1259953556
transform 1 0 1315 0 1 0
box -2 0 476 513
use blankpad  blankpad_25
timestamp 1259953556
transform 1 0 1789 0 1 0
box -2 0 476 513
use blankpad  blankpad_24
timestamp 1259953556
transform 1 0 2263 0 1 0
box -2 0 476 513
use blankpad  blankpad_23
timestamp 1259953556
transform 1 0 2737 0 1 0
box -2 0 476 513
use blankpad  blankpad_22
timestamp 1259953556
transform 1 0 3211 0 1 0
box -2 0 476 513
use blankpad  blankpad_21
timestamp 1259953556
transform 1 0 3685 0 1 0
box -2 0 476 513
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 4487 0 1 367
box 0 2 511 4264
use blankpad  blankpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 367
box -2 0 476 513
use blankpad  blankpad_20
timestamp 1259953556
transform 1 0 4159 0 1 0
box -2 0 476 513
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 5000 513
<< end >>
