* SPICE3 file created from 2-OR.ext - technology: scmos

M1000 a_165_n141# B a_157_n141# Vdd pfet w=1.8u l=0.6u
+ ad=1.62p pd=5.4u as=3.24p ps=7.2u 
M1001 Vdd A a_165_n141# Vdd pfet w=1.8u l=0.6u
+ ad=230.58p pd=285u as=0p ps=0u 
M1002 a_179_n141# a_157_n141# Vdd Vdd pfet w=1.8u l=0.6u
+ ad=3.24p pd=7.2u as=0p ps=0u 
M1003 a_199_n186# a_179_n141# Vdd Vdd pfet w=18u l=0.6u
+ ad=32.4p pd=39.6u as=0p ps=0u 
M1004 Z a_199_n186# Vdd Vdd pfet w=18u l=0.6u
+ ad=162p pd=198u as=0p ps=0u 
M1005 Vdd a_199_n186# Z Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1006 Z a_199_n186# Vdd Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1007 Vdd a_199_n186# Z Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1008 Z a_199_n186# Vdd Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1009 Vdd a_199_n186# Z Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1010 Z a_199_n186# Vdd Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1011 Vdd a_199_n186# Z Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1012 Z a_199_n186# Vdd Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1013 Vdd a_199_n186# Z Vdd pfet w=18u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1014 a_157_n141# B Gnd Gnd nfet w=1.8u l=0.6u
+ ad=3.24p pd=7.2u as=119.88p ps=165.6u 
M1015 Gnd A a_157_n141# Gnd nfet w=1.8u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1016 a_179_n141# a_157_n141# Gnd Gnd nfet w=1.8u l=0.6u
+ ad=3.24p pd=7.2u as=0p ps=0u 
M1017 a_199_n186# a_179_n141# Gnd Gnd nfet w=9u l=0.6u
+ ad=16.2p pd=21.6u as=0p ps=0u 
M1018 Z a_199_n186# Gnd Gnd nfet w=9u l=0.6u
+ ad=81p pd=108u as=0p ps=0u 
M1019 Gnd a_199_n186# Z Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1020 Z a_199_n186# Gnd Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1021 Gnd a_199_n186# Z Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1022 Z a_199_n186# Gnd Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1023 Gnd a_199_n186# Z Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1024 Z a_199_n186# Gnd Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1025 Gnd a_199_n186# Z Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1026 Z a_199_n186# Gnd Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1027 Gnd a_199_n186# Z Gnd nfet w=9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
